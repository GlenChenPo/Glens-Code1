`define CYCLE_TIME      5.6
`define SEED_NUMBER     321
`define PATTERN_NUMBER 100

module PATTERN(
     //Output Port
    clk,
    rst_n,
    in_valid,
    in_valid2,
    matrix_size,
    matrix,
    matrix_idx,
    mode,

    //Input Port
    out_valid,
    out_value
    );


`protected
^Y+<GC-K4DM.Q&31G^aTW9GEG.A#g,M70I-OKfL>g29[;[Wg14CG0)8[(I.T25?3
gI):d&+B4[NLCPecJea??JY<@S5HV[H]OfARZ&/7fLTbaQK3HCKUd^<)90Hb]DP_
dFe5<D,QZ3A<+-gX8,\PFC]99LMFIWg-MeUJ[^=SBT5MdT<JeJ)9g^=\^K_9CWVB
4DI@01&+PbN,F^JFdRI3#SJN?e&;<<g&PJdMY7QS^M3VV0&+b5XZM#F)6f;:QA_V
C6PA2-)Z3bRgX&a.^L]E&_H\(:E^X1^.U-[cNM+2^;XVH$
`endprotected
output          clk, rst_n, in_valid, in_valid2;
output  [ 7:0]  matrix;
output reg      mode;
output reg [ 1:0]  matrix_size;
output reg [ 3:0]  matrix_idx;
input           out_valid;
input           out_value;


`protected
O;^#&R\,=e38E@g[,V20(N].J?0<,gGM@Y(RIE4)LP)RNVObc#_+-)GeQ@5.IHZc
\ZfRUQQ+?F>6&Y6OWWLJ[K8c@-ZP>2^38>)gVA:f97<.DbAQfZEV4=WO5ZH219O<
S+V:D#4P>R\]R,H7:[\-,)[:4+N6ZOJ(L\2<B_b83#3EVE&c\D]3B,3QfIb1G7[]
O7;UX)G8@:b+?8=K9.FR^^]f8T(?48b4Z+4N<&-9E&@T=4bU_VHC1##JZ[X8g?1I
&&@K((I],#KQ+/&=B=ccJ;Wgb[8/)Z]HU<#L0LDYV&b?/^D#>L1/Z@9R:aFRRRZV
R86@Z;O(KeU,<+RI)]6QA[>NC\=&F_8BLe7Z0fE0fHX;+JF^&62Z7I(V#BKIXRBc
#_I,gH3U92WFGf05#LgQKe7Q12)Kbe,7:SZ>^4=.:#+J[EI30S2O<?ZfFZMULUW9
G=B>Q4Pg^L?[6S6T.0WGLeB#L_R7+A##Jb>XHR^Ta2^[M1)9_3,2[4.#9aQ#T>bA
WN23H7O?Y0QHCDga8LOGTTD,9BB6]bXJa;3aUM>&LBG6QV5;3,PFV+b+,(6\<b<A
6BN@O=R=d1UJEKT:6VLEf-3/IMfBNGfF_gZ2F?45^@T=(S8EI6^JMM_@Ge3,c3S<
P^1_NEL?8OMQ>-ff_0a72)AMEc0\,X(-6(M]VS-^B)B;F/8?aJP-0[f^,E-8#\H>
)=DW.R]XL=P9H<SJB6RI=AS<WA&QWX,beaZ2N1:3<\VV?9eg#<K(]d5JG[ee/+C.
d:=>CHJVM1S(D5D;0L05;^26=UADbE#Z\)4+J?3g(<Z.PeIQ=REOVeGTbY>6CXT?
TT/43&[(OSCQZ<;dWWM5g<]EG=-4e#&Vf7>/8RXXX^BYUF-Le4a.7VJ:C[XfK.^W
Y&I5HS@g<O<[?3PT&X?+W+1BS-2QC^1ae^&Z.9EMPFPf\ea]bJ[#TC>bC.,,(ZHK
POF\OfX[\2#b=A6Sg4a^,;GI0gSD+S^7=8ceY.S,Ac+8<C=K5;4d4?DWB(d>UGTB
f@_KeccP:]+)PZ55gFU9a#,;\1>Pf;Ta6>^]Q#f=;-VbGK^FFRL>,1XdK(-L6&\M
#_HGUN:1XB]_-N\)BPd[a8OL,[1J^WgT[>^GYZVYP^&&3/5G.9Q.EC618ABKb:Nb
3D&Q=DY9)M[A\Be6E-a_P7COB]9EKZ\8:L[89H_/FF0DE,?=H3Y;-X^CF/V]bd.-
LR#M+6RG_\/FfGf5#f6>9bJ#GMXN9b&,LN3]IbN;)BDY,K93afa/P+AS&SYLR;I1
@=_BMPB:JLD-YF8XD9,7;&M=7?B3&)Z0)AR#+2eST4(Q;H;EWMC8?PgJ]\VRTR3L
ZZ>;Ac=3Y_1_KAc2:RDZ4ANc<a,FBVbb2Qa5^\F?f7WeGGUM<68F@_9[[B/3\/bf
L:bWM>JA(FF>\,DM,UV:C9_GfaL?I\[/Pg>@L/5c_LIa19J^Q4(fMR+?_OL((_Wc
c]H=D?ZT<))#/EF<O&2.S:Q?.bQJ_Q89U/N</[KL<]JVWL=fIG6.AFLE(gG)XP4X
f>_QgV/]8#>b\BIPb5d>#L(7aOR[d9bd(UH:]BI/Z]1&Z=)<(6IHYDANIT)UDK(E
G[^&=1R1PZ8S#fM+X5#=Q:c,\FfL?@eV3/H+-0KP8(Y6;#e:T+[ODI,T)QPFP6B,
7dGaS5,UPD]6\1-D-;/FJ/W7^1#0-RIad[;[GBO;gYA0DTHZ_])#T::DZLMV]]S+
54bBWH)0GNE8H@@9dR^1aEc:G/E.\,LRC4OJ:Qf^WFgZf?SULTJZ^GIfX[NA&F?Q
([J/g2J?1K20/Z0995Te)@dL>6P0LQ\QId+c]bNbA@Wd]/+-Z@OM(gV9>KIE8U1Q
@,G(.#c,9bZWBS=C1STTaL1VSC/c16]cR]AGBRD>3<3N=WEg-Hd]-3IHOHIU:9&H
Ga9/BXTQWU<Ja#c#Z>6f.O)X/.E4.:JFM[Q1JV5bZ,SVHLa#?C6L#=Z],^\cWO>]
68O[4d4NDLWBb,8eH\<6>S\ZA2656GGP_cZe7C/AFYce,IWEV5(D12/1MIS4W>C#
Q-AQAH6KRG>bRa/,,&+N&)]]:ZSZbN9](#F17<OVG(+N95#F&:ADOgBgAX=X>4)N
SLKU4UJ-6@WB&9_<cSZC;>#=:4I?C1aC6ED^_=58Ad+(g@R8:E[3XUPQaB&W1Db9
O83cEI\Y@+fd0T:;01-]eB&7aBPf2&Z0e86ETcYF0cAg;H&VAOL6N5O4g62FaC=P
Zd35R_@J^e-9Q7M6)>L9E53-,<HG8478YDF\O8eXI)0I??TcS:b7-1LK2KBAcg6@
d3dFXD\,-(E#e,:?X]Db1BAYJ<O1fFGA_CL-J)LScO@4MeB8\bB<+RGV9B@8+@7#
fLZe(f\BL=OZD8M4N]]C++Q/WG&_+ZgLa?TX^GTE00G+cb.40,fJ9c)A;2Pd@OGD
<\VG;>\b6;G<YTY=b(bTN;>D9&5[^aNea4FB[a)-gMeRg2Y&_5,L]fL9ge70X?UC
)IS[+4a44O^bga6RN>/)LX-E76#_L=)W+E[\3<d<VZXB6]8e3XQMdT^b:B>)(aF5
GFZXD:g&N_MHIMJG612@O5e84F,=;#>59:)MOb1KDL:^\)gM#_96^YVKCJZYM^.3
,Ab+?^R0/fRSQ9ZK6HFCZb-8V+-&=]YNfXCEEXU/N\6-[Rf-bd1GJ3NeC&NOYHeP
1S6X[_(U(>T0-EWZY,1>ZL<^cSe>MPHGOR)WLMJ[UbH6RU>@da3c4Bef2>b?Y.CQ
Va8?SB<6VNbYR::1RO;R8N&<H\U<)C&8TeFQJTQ+P(.1g)/(N=<^SB)@5e;(&WE_
VNP=5Kef<4<SREX^>;,V(a8D=?39RaA@<6]3:b8b@[C.4_Q(1C7(:Sa,88>J;3YK
@@b)e91(A,L<=-L+;#^+L/-.PZ9+GN--?HAN;LY\#7;g05bd,SNRcY9G^TNJOOdI
IM^7e(F#O1O0(U7VC>/WXH5Be(deSd,ggW&E@SZJ[(PT+L@F]BVB:Yb0507IHC&.
[[)7^WA_+KQ4b[Id(PSZS^MUXWFMP2VZ/b-FWS-F;IQKgAdW]CcRJNZ)OYdJ&@bJ
gBD2DgcAW<?B&>+3eVKJ<dX@Qd&Z5?(cdGb.\+b15gB+4L]b+XL-@B:Yg4Ia#KAR
Z5bISIfECZAA(RX#T;@0dOE@_FYHRcd\5QKUKVGP&,HM^AOR_)T:^eS^WXQ5OF<d
0\(]/CRKCg>P#;CDc<48TKg8(UGK<3g.2340E2bgg7O^:08cGSW#<McH3[:D14a(
)_=PLW+P<eXL6CJ7ZFb\dX5UYK>\0e#>d3@)\&_HDRYK;R7=JS>(MP9_S=FYY@Z+
J,4/1([(S+,&6.U5]:QIUO4AUCHF^e#/_VKDKdc&,K=Xaa8-AKF9:X<4W#3=W6P^
K]+D];,IN0Ca5328P&8H7,BQ7C-29e5eP@6PG[N.YCPJ9K-B-U-5;H3d;(c(da(W
N^D3)?O-0YNQX^F.(9I[B<FV-1T4K[I]BTG#MCMOIF71&f6d8[1]\K#Jb^)/,eAR
V36&4<D7FL[CD.-_.DVW,-UA3>@EN&D/(K@e]CafYW?V<G-NLJD8c2>HVd#/N]\(
Z:XM1ZPTFC/UL.M=G&fbBM.B<O;WBBW>S3J4X[N(#?0,W^#Y0O4BQcS9GLP&c)6b
IMK8@6B5OEgB&GP,,N>D8@c3_gfd.J1)KTS9gL98GJ8(B(?_)IZWc.+Ec#)S/:Y+
X9>@:cO^XTS0b><T4:F#.a0)e8JL=OKMbF>:V#JXI[HeH(-b>gX.dTbZU<&69U3/
N8LA582c<SFUgA3_daTVf_D_ED2N@;J6]Xbe,e(.Q5dE8cJfPNR]U+(S@If@MTG<
b&<C9W?A59=P)J)SD-B4a1c4=a8QD<35>>G[cKgS6a<:Qa50:+RV#7S5C4O^gA4;
VFOP4]]8OMKcW9,5I>F0d)_UcX9G[:dJ6[N489M/T;C@/c2DAdeW]I&KY>@.YaeF
\^N]38>HL?b=aQ1Lga0gafZd2C:)IJQU4N:_IC^+f3+0Y_U.#&P]4PK9AAIS_^BN
7@DTGW-UI6QN\Jb.C/YB(OIE-=?YH&PKNI+4FeRK[<HX8B6I+JJ3]]X7dfTe;RBc
AaRD5)=.aDJI^25@G//0X@?;8@N+_FgI?,LFg.M;<@26dRTN1?7AO_e,])T?:S#Z
[X57L-HA570e>5=f-\b8]XZ0,->F2P+M1Zf;YAM=W0;eb_Y/#&>>d:^LB=F(XBXO
?[WD#_AU:#d&PWe?JG:S_7@eE9D&-A5IS38;OTEKRCT7WMHGVaWR3[C0D)#Y)c>K
<RBCZ/P58M9=RX8J-X#N6)#SH]Y5G-<M9Kf/],a9I=2P^LSREQ:]_DUP3PJ(g<R8
LU^W03\H8,B;BOV#I,7eRe,>2#5<O6<BYZGA];:#RFf9W?Z._=OANB>;WS-94g1H
=TdU,#dC19HEH<&Ved7)R7YU8e)2M1+Y/@8=-NC(@/.XG5\.W-e/ZOff84W)5Pe1
2PCS9F5J=[+E^T+D\_/E-[A(V?A2L>)bCg](5[/+[2.1ZZ4KgSG_R+Qd-7OT.)QK
L4,94@V&/QIP75I0>7MgaW>&V0XM7O._#bS+1P9W&_^KFZ[,d;/e5)@9YD;)H^#,
Mf46NS2g2F20Vbd[K)cecUA&^:J8E8f57.UZ;XQ9DY[NZ;HfG]>>O9TS&0TQ2?<)
5OPS_K4WW)W-\IU62ScaT#GXa^Ob=9V69,/#A]a6-#L&]0&a35;#DcOBF)(_JH91
&XK/GCEGBTGbQR20=-)<+@E\[HPELJRH-H+MJ@,)Y^^LN)#W[(PG&RcV/>5KL??L
Pa,eW#.=Jde?G=YfF?YQ]dJ;YdVe^3c,gVXf8XN.#>c+WKH((a<g=Q-Q^c1PfRNS
OQ#UVQeB1-a]96.UM5E:P1\>:RXJE3F1T.8c[baJCKM14f15XHGVR]I97OW2d&U1
[7KaKb)Pa;&@;;Ze\D:SKLLJfND7D5Hd]Ad:HAO4RbP5R@63IcJ?MMf^4;>9W-O)
5J-&LVA8[&MG\W,ZVZ.0g+VL/fAS:3T/ePMP.?BcOc/\SZWA:YTVgD(_K(F#V+Z3
L2RgQgO/XUE?d]FLbK:)SKMELf66[L(]a[FJB&Y?PI,#/5cN@0Q.1Qg+,&T@B[;a
EQ8O,MWB455Q\QM4g\JZOR3Z6eNPKBL#0+)7ZW-B0PJbdSO=b/-^Y:g<WDP?.bJE
R+ITNbFgTKXAgNADAB20>7bb?e43HY\KVJY#4Wf]IT1?<(R+;[EO:g+S.d;25I[\
FdO?5.5a:GY8PDfQNS>XD,5HaER=,SdQ(Q9KR@=E^EgI]]#Q:D^&>J>cKG0fU\I<
M#8FBU_#g;45S_X=OA3Q^L48Ea^9JRV15,]+/GBa@1_2>/bJQM:_.:cOd/]&+gKG
6CeXRV;e5eW\fGR3J(bGCcX(ENF&UBf_9ZZ(]\3)+H,TN_c&Qc#2\+KeR/[F7eVF
a?RSdPd#g==Y)KY#5Y/9HBA7GM0f#fdT=4J)b]F.VdRDQQ]<Sf6f3QS:ZA8/<DG@
F[a55.C\fcaIK+<9PNY29K5=J\-EE1961?G;HXOIF?&gRHY0cYE.XHUe2bbC>4XR
5EXg[0NJ)#W:3ICR[:YQ[)^I,)ATHA3#&^F97=@-2@.9a[9;LY\=HBE&+GePRT^<
FaeM;5e:(Bag]:-3a>V4UeBSN9aUGDZ#V?-Z(E9fTSU^,[@PK5I0ASO^a7=38.<X
de[Y2_.CSf(MTHJ2O=@SUJ0;+bXMbSK>R/PbI.?U;Cag\<(U(eU-<GEA]L^X5e^=
JF(AA/I3/D+U-f\11a0SV@:=gY5^]bc.G6cR(RO.)eE7Y<D,&FSH==-D,-DFO/K)
Yg3Q.58c3bH2Id=1&eFG,fVG=bc@_8e[0Y,Gf&F.RI-C>?[R6\.C(4JTe1:M/U1W
M3H=,@)XFM6T.S+>=VD9:B<O@0B./IVDH=XKAM>O[c-gV.c?QHO,B6Y@V82#]),5
IZ](&1D;QUSRFKD3-@-Ec@B>F\;YL3S6/I/V<<e>AV]/Yc^5[bW[@7K(AJA2/PH(
CK.I70:L=,_.UL-^2Je(V?FfHfIcdQ6EB>S]Id=2U,eQL7K._][^R;eGV1WSL+DK
5cH?2P^CIA7<;)R<g2Qe[GP((?,a=41B8PV>7Q8ec#-L-K;,J&4O?5AL2\S1UZbC
X0GAIPU/>\MA<?d3dJ^0?10MRT9AE+8-c5^[2TNf7\YeQ#U:>d;&)IOH;SW-/g5F
2FbfZJd(d;N)K05a^Ng2b>&J&\#]-80c_RR9&OHZA0\)H-aeISAUP/@S1?7:ba]a
_RA5PD_b<-KaL>#>1ZZ5eaAag6XY^:B[I@ND=1gb4?Ub;73<e++9f1aU<JfU2>\G
fW+f6AK4b6H]\Z22cYa3N;C<^>D^]XP]XTDSgcG;ae\J+U<BFBeHcGI87GV<?[BJ
f8MYaPYcF;REVRg2ZOEffB-6I@,Vf0;),R>5PLX#/K>I;=/&)S&-7OK3CcYGD97g
<;7CRHg>aEa+6P#7.bFELg+Z(g6HT&Kcd8U12g=d7\M?#48eeG=]I;=B<UMf6A4>
4R9G.V@bPD2=H,LF<;8W8AYBQQfY[T/8L<bT^T,g^Zb5OMaE)\FeaMAOcfgL]>M5
EN:YL8)M\\;6M-@aNcSQ,&CDBKB\P/=KK5TBY7Sc>-TVAX)T5)1S9^SAU_fW9cO=
;26M\4=G:O,<Jd\9eX,[[cZ6F476-.IdI,>XZ,,IA9Ba0@;3M+]f.]#g?f@&&)Ue
?gZWV5@#4eNc-)L+=OfMQ-a+_RJB^XFT592_T(aL+f1+U[f9Je/D@Wd+bGTN85R^
,3G][e<8T&RI[ccHTSVKJeG4VBMBYH+2:<1K8.;47B((bd[PU-HQZGQ2]4N@-D:Z
R2gR.,1,:b0N:;W?N<5--?S)f8>0?I,G[GI#Z7H8dBH5Ld-P@T.)\&5ceM/(]3gR
+;?d>\@#cb,F:?Z0BaC<<>/>ZU-TM<X<ZCLR>C74DN8<0=L65ZNf1/N)D0Z<^RU0
(ZK:UA=8^<UI2^b[/<\0Id@,02+d[TbZ2Z01]eXSdUKSFU]MJg?KO:@-02.L+=(U
b?OV#a2O;+JBHeOQaa4Ea6B0A^9acLb&Wg]KVY.=BMUTDF.cSI2KYS13bP@85X=>
abE:.VA6/2Z^IKF=^DW[IXLWTY0Q=\V>1d#IB@UfI]eJ?^?9L?)[\b=&U2O&PId2
)W4g(1NWY_Rg)b<9ISf@=>[TR4XaT71f?>J/GRf9GO:0d;)aKVH>C0IfX78cE[;;
T5fFW@03Q+(2,NOa&<CWX,;aZM\W;^f11)Y;FHIZ-U4O+UGP)P(M&T;:LF@N.c5,
EMN(,0e4T;PRF4]O7b[:<(?3HY44NKL&8O,R^A#+2UI:fNeJ,OA]DYdeRQ^I#]O)
eeNE4@P;:+B+T^c7&K+<\))\7cP/G>@+Kf=dH#aca7XC[@/C)>K@Z6<,4U1b1&#g
g.LJE+NNA<d;YT?&M?-#0/-=_QI+RdeQ_9[1,b^,CH<1-D=FP0P7gJY(dVT=MZR@
ETce5AfIgDBE:F#bS;T[P6eLGHYM@A_T^W3KNFS2@6>9#a0WWQ^TW\?b)FDa=W+(
U_O(T+F\b_R/TC42<^M@M:XaCJW[6Q[4cA8>O:X<+25f_T[,:6E.OFJf:N(Zd(DK
HW,0bAVg@=K:]YM4WFGHVW=R[1&We?CW3O/\GafY2MgTT_VNY,)20#36<2>>YD<&
.29ETf5\>XAd_GAcgC,2L_4?(b6B1Z;OYLMJI\9,3W;g8MI95aY@GM,56#L(SCNK
a>#DOE&)BV4?(30<W3-6bQbYFB_KTHP@3fW9Z#=DOU6EK?>O?R36_R/>T:?7?>^<
N8PUS9[afg_AYK=MH25_M0I5XY;F6E-/JT&\7G5_W-aBBU[XN-a(68:35L]?d4G<
a_C\5+4V^DM/G+NT)H\8HWYQJ0;ACPD4^C>U^P-?P8@RDeLAc-<U+TNP>GL-<CDJ
M)-C-G[VEg+.bBbSG_I02H0#)1+ST&bJeK#,[PcK-9a:3fLB&@c&5923HV##Ve=\
/U_dZ7&&W7\-gH,H+;X_GOY1AE/#1cV5,5VYFWD6.PNf(6PUQ]35UZTM7]8[634B
+c58=c7MaP>0]eg3NH]0B<1#OL8f2>-UE)@GHfT;@\IAJd<1WgK;:7J_?K\LbH1/
HSG+?.7<:[<T2Z]26=(>EfJN6g-N00.C8-;U),7DVM2cc=O#1dfHed9aDC@8b.Qc
6dGf=.[G9YZP-:+P:@24dfUdfZLVHJ:f/M.cFN<H9X,DZWZgT=DXQ7E^CL<Nc=dP
WBXBJGD8S^=ZPBC,O_:dYYI]&:>L#U4RF5S40T=:=\UWL+,PBG1@^@D3NND.9RL^
]?LI/K3Z_WTdB9Ve2.0K0SUG&Z0QId?Q;)M5=1U/UX.KG2)F]0&#gW7806C(FZZO
[;SQd[T((&Dg>3,)TSA?Y^)1IEC/&,JCg664+D2-E<6g.M;<DXYN,?bNGP,J2g7\
FL6>=S5H7c;@Dd7NU1151YbI#<4B)BGMZ7MWP)>&.T,NfRQA1,eg]5?bV+.adS+e
C,[P2QS1+:VZPe^.Z2YQfG6/;DD1C71(+9RMMZd3^4[aNNT23X\51e[eJ3+Iea6Q
9EB7MH)[CGZ?VfBR0>+YH^GJ/)/EXL)KgH@AI,9EKXBW?[MA#Ob=&_\;3^HM4^g4
dHP/78)744cO^QbTbV-9&8GXN]A1Va.&R&#b#8(e\/UKN:KW3^==[4PPCU^9GJ#I
f5f?\C5Mg>5d-_AHTd=_KLA05S2:C_aK6UG@9?Q@HBC3gVd_M\d4cb<>Lc.b=a9W
__K7NL7d1BScNYL6E_\dPV&bC4N8fHE9C_Qf@)<6L\Qb,Rd+N\?0EH&/6=MTYK=a
WMMYC/Y<>U<#cEL,(2P?UYcU8(&dEB75K>X-[SKcGA307>(e.)83OWUKFRHLADXb
O4S;Wd9Id/Kcg:E2J_)CAJ>:E&9bMI?8/bY6NK=F.B.W@LN/8L(Z(d_7FR75:X?#
F<[<-I0C9FY4E^SfY,1X+J,f[BLJ+WBH&IEF282#Q6d@3I1&fE6#cI=XaFM[@JFd
+P&Qa0H7W[3?QfZ6>-&=eP]7a(:Y_\R@2<GQ5BR<:L^Xea<?M>,^<Nc4SQVCS75#
B?QGE;A=PG<K7P.>8YR(RQKB1H;-E^ARa,\0\DbJ1ddY?gS[(T#2UCN\dU:T4bTW
K3N/,0FSfT,6A70a(:<WO@XK/J;@DS5TdJ0H9F09QY@^9LI:)@+],e,HbEdgT7;R
[[RQGa]Md0?)@)XZH=#UPbUU.-48OZ[K>JY\R7_NMdA[W1,T,A&)T7^]?/BUJ-,U
;V7OY\Zb_DGFRb.(>4&B/N>@dUL6f>H?Me;FOHPb\@g:CZc3IN6D8INSQdcW>2:N
:UCE)0-VN^X.f0E.#ec5CdUZ;\=2]#:NWc#;GX=IG/[\-=(=L^Xb14>#QO69F,FL
+C3EGa>.Q;DEGJT^;VGTB2b=P3)^C(fgTXF<<31U]6g):GeYfDK[#G3?7H1Q+<_)
[FX+A)8&F[\C:IH)#XKR@MSZ:NG@[^DWY;4eaJdV@GaH(<M^]IRUNZMI<@&<3=U>
J=&P]eKg:IC5aP)YW>I827<G3-83H?OS2#A5cW<C.D\+BVGa/7W7J[Sc:@fE<)X,
]T;ICacQ/X,+N;a]#TY?#7=a@3I\c)O8c4015SWgO>>SB3\Q1\+S++1EE@V01D1?
##KXW58ZMQ2W:O16&]7]04)?2GMec0gTfMWcVZDO(?3CQ(1@OKP8-4V0;4Rd.fQ(
a#SgdT_eR&8+[BV01dKS=.9HNH<>CH^AFO<),J/6.+[_=4C&3XO>SUd&KFUS^+,e
C>VOcC)P[7J+I:(b6M-WdW2WO<gZ:AdQ[V<cdO9KGdJFa09L4WL.OZM+T2I3N9=f
Z9ETPDBVVQ);DF3C9W@=GSGY<f2M6FA1B/ZVXTWGLW/X4bg-b#D>[BQA6R3IANYL
J-241<GR\:f/c3bEE.-+I/@C>RKNF?dfS<?4dS;XPJGgE@ND1J)]S3Ra(TDbYUFG
RE4gJ<T4YDB7DaNaJe[b8f(43C22LfY\^fd-UaZ3W8R>1Z?>9TD[c90AC]fR@7F-
]b0dM<XO?4Y]?W>4U.M>\10d9DDcgUTaM8WUCP.YSX_Y(J^0/dHBAQB+&S+-8VP=
OEg;T=EIDe>456BQ_2Q6@EdCc9[Q/[fg5cd=8/RVEI)6<BU8Z=:A[U]f)+e@-d?(
8;,JEFATb_@;LT0-10<(Y16B/09:FHIRcVI];3PS1RTaVUA)]#<@@ZP5Lbd&DRR[
:ATA?<&QVZ]bFd>B^?/DTbdX>]PL)?Q@]deRI:M4gN9189JLVEK/U?M75(eF:,a7
,-eNHe=4b=]9:<,MQ2<-Cd:E\&GgH-?(?CgK\B#O[Bc]O6f5OPP_)\S6DJY::R0R
Z_OUMgd+?)T0\T.=8I)[K:-NZ4UfAUZ?[>)Qe7NM<RdKOA5Ma,_e[0Q6aeOF>b#^
.@Z7-TUUaU/T89QQ+.TZFf6(4gbKDPOMXRDBaU>cg_YTQc(5QNc??;Q6KQXRbZF0
:1RS13O/]#B:ACU+P/&A:N:&:E750;Y+eAc5J&&3Q+-S^WN@?864cT@+>SNC&LNE
FBX7a#O)?;G,3-CR@-:@1/g<^7KH#B=.UT0b5fRNX3,OV>6T]U61GA>/QEF?_Y_g
Ne=WWT+Y^TG)EL=]dISbc&]FU<QH1]Kb/JI^BeYZb&f6H/7=LFfF;WL?U8fKeb[D
DB6b^3aQQ:82K4_#\F=JY)e--&Y;Jdg)^5W,F)PWeAKa1S]Mfg+SM267@5?VB)FY
L^RJL#16=J^/MN<R/B[S16^?SRR+Nf0bWB)0@C&Q(+gL5T5BO)#bN?X0+6:a:8E\
U,-<c5)<KTK+9T+&.?bA:FO_5KgRd;QbHcTGJ?/(,Y@g2CPEe4P)(^>84bQg+O]Q
H1b/-A;)+RP:dUMHOMA@17?4-&D3+)DNDJ:AOO7E:R>H-<SNbK##&<,9PWe)<J9Y
ceDX(b9S-TeZ23+&_PC9R,-+[c<5A3B7AgEMM&e284>3Vf4-@8A?[+SM/+bSJAEE
\A.15XA^eM\P=VL<gN5S0Jc5Pe[[U8R.]=fV2bc+edDF(ZY@0O+9E]a<9^#50G?E
TMY<\7@D[WY)[_NHZ3J3,.bSF+1T0Ka94&98(FL_L]d&+KOcQ?P60=EX22I<BfeZ
2GDWfARBBLE5Ld.;37=bTNeg4G34aaQ2UO]D^e-L,gc:ZbgB=+Gd.KfJ+[&^GHVe
7#U7H^JR22]4([N)1PJOaW=.5ecN(MUfJ0[Z]fO@D&:.NV3_@/7.]W-&X3):cF]d
(Lf.N?Lc.eAU9-#,e^GTU=e@eG,ENH1gQX<21EMeea+58OIZ_fMXI-VDBFX-Ff-X
Y<fN]O4C4AEDSOX)f#0KV]:8XgX9PV3RP(De4?dK<Z?I\@W#N6GUUZe(_8,H)b>C
:K>-99:PH>I)S[WRXJM)X8AFRQ(eFc:/046ZEC@QFWW7TA3SXM[^gPD/G,Y#8&WG
3_d>df.a.N:8a81FYK[20KKY-3a7;a-X;P9<K@Qb(aT#ZR)gU_Z740@(>UA#3^^5
RdYYG)W:N>3)04#)QKE-5IecWKB2L]L06N^XBK1<S,6,8>dLM=f^+3@T<I=f,A6/
3-/=.05O;(6H=X8)[3URM@+eLY^&H18_c3Wf&7(<=+Y;;/A?;37aZ-+M8&de:YCb
/ODHMD<^.3T.D4AJF/.BS7J+8[?5H-gD]c:3NQe295(1Q/K/1+1UTC5[W@0gTR(T
K2Ab]N^6(PXTG0LdS-ObMHFH]EZ41Cb[\^GECb]=R]>DMb2Q?Bca(Z;^SA(Wf3[e
FL024)V(:?3gFBW+bDc=V=(]CLKbf-JI0>B,d1(#GFOcJ>ZG],U58/?=]]@&(0[B
EF4I+O1<?<:IR&afbAO6@56&FV+6V0B.-]?+6.U+IV/dIedA@62cDE<;(EB>+F_S
3&+D:P]@HeM)S@:N8V<;Faf7+;=O<6N6NTUBa,,efI\2I\D5FEQ:c7)\;-1-Q(f2
;ICU=[BQ?G-V;CT\3J@#GJd>,?]N9#4N:Y<@?:FTJQgNYR1=C]DV7LR#O\-6G&O8
Q+WC4D5c7d85cA/8/dFJ>g&TJP/OGgaE8U.I/BJ3C:^)1fF(NH+6;cR,Y+X@W)(f
U@8Gc[.XHG1X@Y9XJVSgME.fLcD=GP?@U4U>\^<O+C/Lg]44KW2dfecYcN(0:c75
0R>dT;>a[L41I[Fc>HX?#Ed(S@[)IT=O-+6(025;BR4DU(SDL?94U/3B()@&EYH;
1VHX9_RG&TMF6565WQ.W6eII+XO&SC4)b?(+9-;X-_<B_FX.5>56;OV6#?O94G2?
aD(H>KS0g:3aUIX;):U5K=K)?P>XZBHH>b4P=DcWYd]8[NOCIb8+P@dfS[AS/agY
G#^5?KHR_6[9bQ-&0U,&d9OTQ.=R0dYX1H0NP;@;R/()0(Pe@-3b7R@7_[eY[OP,
T\RRI8Jf7X;/EO=gJ0b4<;S\<5Ibg,:10PP;VZ[+NG&(e(C:egT>QKT/E=LIMTeU
OB.aa48+bXV_ZF1cM+Q.?SH\;e0\:4\KCZRZ2LU8f&)gZCS-X]&-3@Ed?E7\1<(8
W392,L6ZL[AgK_N..HKX#YbM,^0.9BBA?Z:Y-R&LI<ZL3;9C#L^C=ED,V[LK[+PO
dT4R:>D&5DD+BOUE4UKW1NNJg2^QQ\XGF&a5fE6;QS_c<L,DdEgb#a<c0OBAc8+M
&NY?+A^T5:U>dHEH;UVLPeTODaYZ@G5KCX/NGc:PW(TMY6RdDM37>fC6@>_cKfM0
Ia=JAFOPP9]B^#cL08Dff,=W_fKV]0ZdXb^cR4[>DJBbN-]fMgS7,eQ^EIgIg,/&
6T[/,2J\W[77U8Q_&&HU0LU46G&FbYHAZ0X[IK^>E^R&]Qd9:aA<.=f62F)&GC6V
gc4e=;J\BbR)d4G+][_0IddY\<B]##9g8[,_JB])51SQb_B>_YGcU(C-TQYKGJa^
.;0[?eJO9fA-d@7=>(EK4HEF?&T]YIf>gP-UGfR=c==4Hb0?a--&c;P_)VABcO^)
(&OTRY;407<ZQP#PbCH)aWa^^[J(REfSSQ^f>VJK>FY/J+g@_C-)8#S1W<DN&B0T
IW#5>.L[CHEOe1Ld?20]H3>AFaU)E[:?I?B-5\Z(5M3YX^WW173aU_aJ)a@9D(.)
]c3(=,[/6@_2?ca_/Y_(PW)C3\e;7]E/0L6U-Y,NYW2eS)ULEAZ^(1Y1bK=WZI-b
KR5c=?-Y9N3OW6a?6,FbJ:X<BBHgH\RX?\^RBL6IHF6-@Xb8KI/Z=7A>e]4cWD;f
J8;L3Rg7d?W]ad^<=30:>dd)-7S/aTMVRPLO\./3Na5MYYg@a@e;P813^4EHM#OH
<Z^#HX_)4N]5)eDNXXHaJ+dH)@[@ZV=I;S@F0++=H+A4^cEF0-G)SZWFTS^.+;>/
LIC7MTN(H;>><Z8fQ1B3\+RIA&2WGD/5ZAB^0RKN?9MMSbT&:(T;BJeZ.c&PUbD>
^d@G=@EgfQGM=F^TI].2>_H\Z7Df-gV;M6FA&@UEUPKcLNbBSc,VSeZ1+CIcc9Q8
E78S:DNe2b[D9MZ2I>-3Q[C?.-^TPTa5ND@1-<\g-a:CPgeS^UR[01d5F_\g:FAF
QW8b=9?(QM_E@^a?YY76].28;L3Y@e?+V+\UAEJIE/4-g-SbIbB;BE#U.CX^7UJI
AWDKL4C]+UAWT=^cMb)ce9PR]W,(3[DI[7WUf[DNAW6d=DY[ZXUH>+YY&T+<H;3E
e7=\H/7R-Fd=c9H5&aRNQ<>H1A)Q6-1SSaYE6D=aU]RD3S;[<GRd1;>?g8M+0-<1
L/ARP@#dbYJYRDfa25]RTd/-O_^a/?eLd;@Z9QF\\]e=43_7N1CbL;?V<6IJE7[G
C,fg+\ML)60I:S.-g8Mc,g0I2e4)fJ,Cg<eH11:@VLQ_/8M:5fM2AD^bJ#bU0]]c
cQDGXf:]DT-,4_E]NL=.:bDP_KFRM_&1[f7Q_UVJ/U)@?48UF5]f37>Z?RC@0ERO
02d6_41f[.PQU=)VFg[_]V(#2[OJQ0g5YV1,=F3&WPN@D.:RXWb>:DRV>UH./BNV
bS1,&<6,]9PZ6+bMT,[+Aa,IRdba?QBCQ[YSd+0f+.Bg3F_RL\83QAgU;K+;=;gb
FZX1/cQE9T@>IH[VD\):6+MCG-VW>CE)P/^J5a>_.b_RKFYGZ./#bC0/2-_9-F0L
F??;K,b5(0F?d=)K_.^e\VW9U1VD.Q83fH\[E1J>D5DN;,aaQT/6P17PJQGG6_1)
.+E=U:CP>91PRWL/5:,-U4__?(<_0/\?R0W_#U>14307R/6O^SeSaa\+YJ@2QJbQ
R@&?I247]J\-B?T\NXPdZVEa3g_P1DPP]=/2:LCCUdB#\_MCAQ3O>,<\?D<:#L++
.-WL_+U>FK.GU&5Pe2-ea?#RT,I_M.@C?f71H+,\.7(Q(6-PJYR&=U]<Z_T>Z@\5
eY0,B)[4G:C@F,^(86[G)4d)\5cX11@Wd&UOfCL\8F+2F=E_C:F80^OEE9b.56]E
(Y?#^H83/ZXdXNI2VIPVDg@WIO>bXWf,XV60MC@g5dOMV/dP\GU\@+#bT=&5PT[V
ECJ]G.NMJbOU?DdEWIK.GTOR9JV)\A&(QJYF;KRRF<5acTDUH8Y[eeB&\L:RafY3
2==#&[-fZTVA\#>BHQ.)^]+W8;_[U,E@dZ[WT+/f37.C1DOBDJ,<dJ+Ib/J&V/bN
cYGC9^<[_O(,?QQW]4P#(cD22IH7QH_\(YFO[FfFJ2N<5[LQI/H@DYF#6D9HfMAN
A6_BSU^AFC87]X8;(-Og2dZcMB4\d#?3PPPd/_6BAaGMF42;&R1Hb0N\&T?Y[Z-=
:X+5a10D-Dd)Hd#T<LA#d72<WF/G1E\\c3D-=]Z#PJ9J86K&B25=L&\4#Sf.P_OR
Q)^&>BTONg9WJM-&0,a1>IJ(@4\\M&Y=62\#cOBFa/]9^6c25U],@B[J(XQPH<>&
^(X1>-@?gE7Q5(><=&L,3^J;YbIgL4E>?3TR8[UT8:g^YfD)_T4>)^0P=7Z(,9.^
cD-4AVPKIFUC7YI+;0)0D2;ODV.aDBP>gZJ[DUM#0DCaIP]bVgaOKP/LfeE]K,S:
]D&GfHebI[K&2&LF3?9LW1:GU[&IgM6]ZVR[EeVZYHK::ZY/@O-B&).XU(eA9?I+
?SK_0L_gT41=3QABAS..]&;1IIPO4ZA8]+dM41.=6ZF(KPHL&@@0H#IHBJ\EJS8Q
WN>GYcf@@<Ub@\Yg=/XNV;:AX@,R:V.G,QQ5&IdXG(TZ(B[[:K3^aJCZW17:Eg=D
JBZa)AZRe\4^cEV&)#[Z6.5][c2gdJ(+RG6,RaIgZDN.6_cfG&E-T3/2./CRQ,Xf
<?\._6ec^(38J7N##dW71Hdc2>^,3G=5\GDU1Q]Y9gV=D49R8(Z&^Z-B=#U>Y2U=
gEg<>BLdWc:^gcgJN0Y2NZ2R/F7WX1L-0,Uc40Q)4IIO28TDfc;;M^6:cW7ED0e)
_^:6CP@,RQaWf6#fYH5::W@CUQD4=4-,)#8J==S<6JPIa2+R:_K#dUHHcF(9EIU#
9(Z-(-KcWKC:Oa37Q)b&O/J=C_ZUYQ=+,108T)RODW0Q1G6<,:<=5Pa_2Zg90eOc
NLc5?>CX4dO7R:(E63ACZ^6KPORBe@\3Bee[?XPYVdGgEb0[;,G2a5cR+A([D5^I
+#5\A.bYW[U[07?;=2We-<:R;-La[+(-I4;1@)LddRQALZ/A0MJ0[dI4+g<GP\eS
JU[adIFQ13gTJ-2cO(R0>fNYYGHA@3G&U7Ea@+0Qdf46Z@^bS>T]1_(6>ZJTB9JQ
NI)1-(V2D>R=8d17E.NO^8WDO@f.+U_5KeVGD1bSMa;eX49d/0,\aFW_6?U6EF@&
ZDc-#aU:[bJU^R[,d2R^3<SFd-^XR\09(/]_#WXE@)ff9NB(Q+9a/ScGfB,<1=]J
G#RY0.OS=F)Ve7@\^eRFEGdT3M3+L32CN<ZEfNN8>c8>04OZFGULgHV+5+-UZ8,a
V:Z+EfI/N)&R=6,JLTNYH2I8@0:L9>]:eY#5IRC1>8KZ_d<OGC4d]/HKRa\C[NWc
aNbX0]e;^[5>f[#&bJL1E(RR,<](DR>HC5Z]Z.K^g\VfT0;&:MP31#b=2O9dcUC9
@_?PK<RE)Q<YCBCJbO@8KY&^B#(Z-ffHXb<GXSP&^C253E<#]OYcVC/:^H@g#JZH
7W_;d--;G9<-<CcS]c3(MH?>_a<4,)SU=(>Y_F+72W@;Lf](^Gg>?1.KcW?=T_W>
N5\F<V9b[<:+W71gY,Da2;^\1PSLU3+KXZfY6&P)]V>5.F8Cb&8TU?3,E98Z@Z2:
+,&;T#_5C\P1][Kaf#ab,90Hd9B^<S>&dL8I4gT(8BG,CbW+9+E=YVc0/+=D4^]F
NK/WX,(1+)0@EF-2=^D/I+MBe.,(ZUUa(CdI\2)a8+2G<2g)JL9c?Mfc=T5/LPNg
T@&f&fH-E6.1IPMC>:(bO--7+fP008XRV[3S8YQYW:B];]Z9[D.>RO)(>b\P.LCS
f\F1f9aH47DXWG1XAWJF#V<)#/:#5f\E3PE--7B(I+6fKbQ\9OE&HG7O>EdNN7,<
,C=U9:89@g5ZX=-6I?>M1VB(WZ8c+ZdDPd-32@Cf5?W6e36[4HH-+#P3J\-N<c1D
3UUS4Zeg9V[B+[W,WdQM&-6a<IXP3K=R:X#>^H:0T\g?bT45T78GdK51K4Q))13@
-cc7VGU#ac<;?]R[E<MGS<_aVJN94AcODIEb9&d/fAI&<MR6EJ==W8F8ce#ZMga1
7Gce_MTNAg-aW55[);=Ne)O>b^-\;UdEC4=1gF?E9=Y;8OEcIF=9USVDT<18<5L(
^(ecYO]SNE]6@S+5YDA/?7[:.4gG_CT+3<UR4/P>\QR<F,0^>@/_\I2NK0?(8Q+B
(E1=SHX>3bOH;QTA>00/YfJ?[fF6U:5)3?.6#P4F0CG,]H6>TTH39W.AOGg;1#/-
d>8DO=]a7\12AU;F+TPTc<bSGD_&Z(6MR18f3(]#\=2SICJ2a#F]WT?FD)U0:Zb?
c:SI-Q@J;a2RU(;M.=Tc9Df_g3L#:V]3JHYc3A^8,D>E6>>6V>W)+4O5=L(;7Y6(
L;NAM)4Z1P92^7bE,I^.OFH30E]42BSPH\_6/=BWK,XG-;^a1+6_20aB5<e?.c.K
@BTR_.0#X80ML^#JB5Sd=3SEJ;5?NJe[.e<YR&N\3YY6?b1K<.[dTX,a>Gd8e7M(
SHZ\QPZE+\((3bY?:RP:OUA@K3VaDMa6C4,eb0R)BV?F^EcSg:P2#<\:F4NP9Nd>
PPY)A5XJ5+9AUb6_c_38;+HP3KW?()-:ZQ<MbG:B.(;Ube5>R^X?c54U.K=2eR7:
_Ya=]I)T\R=9^OFFJK-.ReE;GB_<<P=,M:2+IIF,ED)NI1H?=B&V;2ZHG,YV.>GG
/ENfAQG;T9X(TBNO:;]R+_Ib8b:a@^H=;\ad&1)F=IO0QVE)ea_7_BIMWaNdPM:H
;(ZB[>5\V7d1I[Zg9R1W9A[<.f\FefU8(GPPCXK@/5<#5ANBJNc0C4E/&Q,S<>D)
GB1>17X\^F:c8cMP[W0V:>Pc#_3A8\HB1gf]He&gf+Y7;S2;F_1VA\>XV:(DFPVe
2.^>ZG9Ve#:f:<F>fb4\E\)PX2^dZ\Pa0;QMG+DBf#6WgD+0B1f\=WCH5<#ab?gZ
>E=XA5RUPNG-f80;250QI:M<bNg91D8WebB&6D@@.&WT&0P?E/D]L+ZQd?OJ_=C7
V9]R^aQQA=H)<;1/f1eH-Z>&K:/FSb0K#D=&J0R]gWK][DYc?Lf+].1/aSKI;R]+
E-W0;GM?GLT#N>#RN3JU5V<cV=T@9c.Ib^7&OWHa/+/DAY3FaUVd+PdPC]F=5:0>
UePRH=DH-97H=USUYAFcTG(Y2S9f;_J::\N^B3e5e7@ZYP1CX-eDd7cB(6^G/:Nb
.L(AAa^J9H+JQ[BHaPA/46d/(..O+a<@YDg1Q_4bNVV5N4MS,[H6<5.bF?;Y/=KI
ZgL7b(6&CD)?JS=P@V(d>S5=Q9W/W5S;R1_F>>eQ@AR2:=4NTdZEf1OCW:T?M.:H
JWZH+_Xg]3@c3DbFd,4[R#bBY[:B2Cc-,XN:Me4+;ZY@IS65)^]N3)]H:+P[S-28
D#7NRP9XY/@)<T&6IWO27G8d+Ng<:>1T6?>J<@eI]0]&^1X.J,&K29FS#67X5\OI
X&[EQ^J&6CabfU@bfdV\.3g;Q+J4):-T\V+VeRJb_<XZ[4@</@J<fA_C(I<Bg3LL
H,1eKYMVN@^UOA(Pb2]#-:UEA@50Q=Y\,_G/RB^f:P>e),EfXf2HcT_3TD8-KcC2
g;/3;=CEU]@CY<^b7?0/V#a?KH(-M7cAHW.)M@-[Z:V=+BdM51Y32/V@]<AfDW;d
Xc3/W34a)Mg&MH#GX[LXBf3_g:/NT4KeMK4[[9KIL=1=2/JWeO#SHZQ6[#YGc0Rc
T@ZPYO&S.6@aLNIf&[R1?N=g367cXUKT2V7Q.8:TXDUS9db<IG3g&C>85cK2.2G.
?fHc&#F1UeJ6I)GZ1AQ#QR,;/.Za^/9ea.ga@Y[R&d=<d>\\S6Lb=&7P&\0d-_d:
1JZb(]3>1?R.,9+EbKKg#N)O]O@JZ7Z5g#&J5H3E\fN4N^RE0A^D,d>;JV..)aIZ
MEU@RC9+BSKFLe;,-g1TQ?DP1A+A/5WJ/QQ[W5g]\V\E/OJ;YQb63_I:>^RF&6g2
d<:T7MOI=Bg58SH?VJ.-GK9(H8U9?52=CPTL_-/<F<8O5e)/J2Fgag24:T4[O7cC
7S61&3)XJ4\eFNP@4g.SbVLCbfdV)Q90gN,;CZ7d6ZO-8N?LeD\@c,UF<)?F2dc5
DgY:):\ATYO.9g5^f1)ORb3RQ?\IJ7=TFY2ee@[72]UP4?8ULZF/(5)fJ<f,9]OI
KfNIW[NW5RB;R#I:XA;M[JO13dL6bCBc<ce1DNA(H47-8?((DRILTEG[;.PIO#e>
(KFc;A,G,TLH27>N_>ZgPN-S_+Y<6-;f]b;2KS9MNFDPO)Z&[DdaB7)HL?dYI6Y1
DLWcABH=;];gg^aJfF_(R9>1:[:>V3-3K^.R5GZW5US=N:E:aWF:D46#5OO)>^/K
X1DH#U#;UdC^]REeHZ&KW;;bK>J)14>5<FeQ^_3:0,Cb0b,5IXH1DQ^7f#.J,\QX
:7=QO=J=d@6W6M9I,:IH=T:6QY7]:7QcfdR;K7:K]O=Z[Q#P0W-PJ,VLCHX0>:4X
D^b6[>)-fY]1C@G4>,:Z&CdA85][)3/^fa+Ogcf-GK+g^PAW]TAbcLbT<.=M[#&Q
&HD0VM\O&:]R&J4EQB8+)#..=R+5912:5a1eDb8Y3a+=TJ;EF24S6+R>eV.JUJMR
IS-#75U?g28Z8UCTL>]7:(QR(/)T16X&ZgbV:&Q,@/TUG3R:?JTN_V2=>88RF[6c
;KTWKgI@dHgJ2B0d3]_T1=E^\d<1d&:K2Ga2UXMWH]AO(M9..X2QR53?0((Cfc[A
c7XB\U<PX+Y@342a?92f33M4L_G,g)-_]b<P\dA<S?R^1=\;5KgX<P?e]P)9G[/>
K(<MB,.+N]e\E-gVG2MAM@_\AF^RYU+[NYCFFN/U_a8JR\:L[\A_NdQQ=2^+\LJA
.H9Qb5Y6L+D6&ESPB40W#J1UMTZ9/R)L0g/fWZIC8TbR8Cg[MDR\IF;FLY@R>V>Z
g<?6F_:Y5RWG?58>NM]NcGVa]52H]K)/\=;3[E]e1#8cB[9A-^XaX;[DYFY;&b#1
B,9BLga[b;S.YQ[BW#>Y6)F6F1#.,fT,V.L-/,J:(80=7Pgf)^XNc5DNSZ.I/G#B
H6aLVYOP+N60<9V;+ag4d.3;d.0fd5ed[[;Q=9E.MCdA-)d;2[_LN6(?O3&ZD:Q@
NM]G9/H0=+.^T8HPaJFD\Z5^K(V[H,ZcQdI:4;^#(=39+NXS[@VSFc[11aa0+Hd<
19?IQIDgJR@bQI\S:a2US5O>;4J,A,8S&9WY/MKEHE(7=;UgL(@+29>6g;_6JgF9
V,>YaT#Y7>;#OC4.2?GQPJ6_FX_\0HF/V(63A\1@VP85C)JLaB2g-?H?UQ>-^Ge^
N]).b)H_QP0VIB2714\+YgTA2@;)(gHVE/VCFJ^6/FS8A(&8YG.M(N,;>,/fY^fH
)7X8ZRaP];c\@+5[(DM88YC,3#HZ3G-(&SD?]?5;[#.X5<M+KJFde5WW/P^decK7
O_J01TGQ_Yd#;?.A&Kg:MV4IWbA7GNbe\Z,6eFSBeU=I??aNU5MYgLeNGHT]ba&b
16Q.YYTF6\Z.YB#-/ae:f]F(UKJQIC7-Md<<BU4JUd>&A\PNG:MCTaM]c(-LF+[?
+>4,;UfAE9REN]1L:]Y;V\9BFP?,B[;3:df)f]XY>XT(9#Y@_6=2NZb;:>aP;_Sd
/_VOQPGG2B1_G1f;4&;163Rd74Jad=DU(1=e2>(2&BNGYE6/QK9U>-FF)_1<dLbS
b;J5G+TJCB9/7=a_)QY#BY&bM7#@Q0O2XQ1I:OI<6D,VZ02_7F./Z,(EMESOE,V:
F??,B[Q<Z_d6<a&ce@GPgX3#1LC@J2>g&5@+^>c,a<D7_fZSLC&>6[3OU+>W6?CS
^)AI(d\EfIDe)+/(KKX[gXeb)a:d;^6K.ceF8B9^2]LW2?CbW-BLV5VJ-2O)31+P
4G4P)0]bL&;FU7[,#C1<3]SJJ>_MeZdF7\La6GDa6R2Q>TOXU+@9UY1Hd4W4^C2F
W2XLde+,J-?YDXYKgH2aE9d]&g286R29H>#<=</ZYC=?+XB+<bF;RQ>T<,2)#]/X
^>[SJZQdOcTF1:3eA@Q+N>@W[&[P)ANJBTC5=(TNYOL7X@d[P5dF_b;L&Q;06_8]
YA41Y[<RBV62^bT6.ga>A8Z_J;KL_Fea):Vd6#J/V_RSbEH93A3^PW,@2QT9S19Z
\Kaf?1C\;&6]KSTN,D1Q1<f>@46Na&PS^(HfT_RA8:WJGg==,7);Kbe[RNgY0K+;
_d-\])O?40X&K4)S_)G#ZVE8b3<8;E2#2^AD2\OZZ&P;70<)HfT[4;e/A,)>+X)K
K+RR:]PAJMJ/&NCZS]cf?FXdZ-+dX^<aB?Y&3Y:7V9d=:&PH.E,OO/;=79MP5U:&
P\]cEfJ3K^,T\N>(@McGcG9Y=ScQGO/CJ)Q?Ta-F<NbJ@Ka>8f/?Ab@F2X(_MF0b
YH>3gAR6[64LZ(,UNL.X4YINH.([I[<]O6ZSD=gBRQ]cIfJ,[J)-MGO3^X7/R&XF
dTe_M8,e,[4=?8PM_0JbeN+JVQDXI9B1=WCR&AJB+T6eO.V2/02YF9O@)F?XG2_^
&/Q_.S?=R.DL^CbCF:CMQK)#B(]G93\^Pc^5OQAW,GE;_GKS#7V>gA@;JEHI-AM#
9OcQKD>-BWEW:Y;\ef^a:MFFaYOOG(HM&;>62\8S^TPY5^#JZFUdY,RWAW7>e-&&
-#L&5MQGQ>8\8<4LcXA2BQWDB(]7L-dBOM)LH]A7HS?b12?M7)Z>.0A3IUX^5)RR
I4[HB9Id4F+M;g8/Y]BEE8,97G=1ScAQZ/A4:a@?Y-29Z]&2&6&bfe2>8/2??,bL
0TUBU]B8FW(8bd1OTdPS=(6aIKb_aQP/ea892I856]WQS6/\b-f6e\DEYC0>?df+
,CYH6AA:F#7X1O5[4._a=Z7\/@@KdEFO5LBABAe/gb[WO(J]+f\b7_&D\9H]E:g.
1+C[CX0T]WLR7K+]YBLD83>b)-H?KM=<.A&0DB4(UG?+9Q7KYHT0Z]b@;P>\T-QW
0<2FT6^/Hc;@:-\>gPW5@Na@6bVe6WI&DL/f(Vd<V[K4Jf:3W3<1.R0a_M0>TYfG
WT(3bR4Q@]a3cBf,@(T;M)dXd8Q#We_,TgZPMdUXM]R,5.?<YF+4gGY?HT=cO?-)
7\09^JO7HK[PYWF<MHfL9L96F=57(@f7edIO/,gL?GN,-U)Fa,+UP0W).IH,4a;/
OGJBBfca3JQ3N02C2gLOa_\AdGN4IX<)CO#:QX)E]8a#K^9]QY^747343RI9QeCI
@9&(&f6CAX:_A_JNS[(BK>I<O_D&J6]d7J:ee]S;ZH9cL5L(D)9@U+d^gV@gC.?/
4CO4+Z[QG)Q?cD?;5#c#CaENLER5(-]P11babC^bb-4@HIKI<4Q@T&Bbef5:>4?&
W0SP/NJdPc1&+,C]?gD>),KB2eP-#aYYFGQQ4=CE9Y_P0;;#eJ]QMK@]>9Z947&Y
1N5aDZEWS#>-YJc6J4>DOY1#6S#W/.P9f&6;QS<D):[70U(VUQ?(IA)3<D39\I-V
)6>26@?,SBZFR+.H2:9NQ-_WF1-,K8(Jc/[9XZ@aJ1Ye_b;8(bVL&eQ8<1KT+]1X
JM&]MTf5/?eK?b@=PDCVQdI^6@eB5&5Ac09;.];2/NY/_^efdXS<:M+?=d\W_BT<
8A@G(9AV55[9@NIbBK=O/Q.2P+E44E=GM@=61cS[DF?-1QFQ3C9DYW+T-@?IS^.d
5e?X8EVH=MOFfdEUT++>f666FM2^CJE8<5(_>fX_=<?R?8@LFOJd=1UH2GZ=AdEQ
F+(I)Q,;Q>7_]5C8.U?-f+)PUG?M;2LZ](/&aJdR1_;KCdfD^F3edVBcUX]+G2+Y
ED@F.(^6WBX#aIX2?4]=gKY]+EO/7g4YJJ1NQ;b.:[AJFL#JXH6184K62KMDP+<5
S+_57:=:-&/gb0[VIQ.NV#N-\7#<XO>W];J=Q4YG_EEGOOPe1XF\4deeBfTIGMfE
J>@IHg<?f./bdC<#b1[R^M=Db/&bH\?>0J)_J?=7/c#e@d+]@1D.9-[R-P:>)B=C
:7<IL=UC].VIZ<BNf9GROTF6MW(gNVUP^5d6G_B<HQH<)BZP.AMPdK<Vc#>KFJ,@
GH-4AM&4+RgIYAaA/4S-C_P2a)/WV6@2;:R\9,WJGRFBYfJgL<CHb<:/0J3+)U:A
,CKZZI020/@3[gg8.f&59+U>M>J@aT:e2JU0AV_(8,IfPHE>G=G)_ZSO^D_X=-@L
//f7&D1-Mf8ZPTV^QZ&^\+7ETGA-#9N[+;OBAUEeS?6+;:Fd(geSUHLb)-.GULG8
a2[b0@G+\0(_1L(L?J7N7gZg;B&eKA;I88C9GL?79@5R)K+.5LXF8@5A<#NIZV9?
HB-b@7#/?;/eDWbRV?/OgO,=D@>KWI@,EDK,ZJLgH^H;I,SgHSX1Z4N:?HT325d+
KX(;0CY2T/WWK@I7LGe^7OPK(4L@W3bH:AR3DHH@_.2Z(dH]FM-)XeNaA8;YOeH6
>EK:DL+RLZf/K6FL3@DPAgG1agEG=MSdH4LWP0e==U2(ER;TLf>A.8GPSYLe8c]\
>QCf03@7T.VHNUAYN^g/@eMQ7cAH+\T<YW?=9Wg_eJ)K3a:g1&V^9G)[&^:96.,I
fA1Q<@@+P)fJB3<6c(EJ&J-+NUEE.+8_N>_adYY(CYRALBa.94_U3UGKRTa1-1Nf
NX2NHJ.FIKfZR<@(5e44T>428>MN1RaUU3;RWTfX5UH64c^8Y@X_CWgI?QK.4#(V
<?JK.Df0E[WdcYed5R;CZ5#.&dTO,9@X[e_-e07]THM2SMVg2A2<E]+]1dPf-CVB
^1T-^O[D.O?;S<+CDSR\6=EBa@+d<S6.,+01<P#WR-I+TF5@(276]02]L@Tc-?IL
<\9UHUDL=[6Q4b2\8?QKMQ(:7IO@.>MP=A@FJ))A8Q](VH,?/ER(T?#IeC=;L+f_
>_D@G?D<>/dL3(6TDOW5SCGBYf+ZZbV(;]UbYU,^G9\,I\V+JTLGS6Yc&6&[1IVJ
U1IFN^&TZ@O/QPAG0F27/[a=[&P#]:=Ldg>^:PJ8EJ25f?/A(+U3D6>]+Z@^]c9Y
^;]0?6cX2/VL1/fKD_#P=A?;4-SA_MdgSd]0G?DBcVe2eEJRALSf#F:6JeeUVf&N
T@\^&I=-.:.1,2^We9_3<-RgI4aDT8BX[IK7/B8T2+6\eD?QTQL3<QDS4EfW+gD4
1Ge+X@2_RO(da.g.]6Z9-68HMDC48c+.M65ZJ#4&&f.._\gb7\C<W-Z2VIB,G?YS
=R-0J;W?=XQ6&F-XOQXN_CO?c05<LC]@0]?9<^WI+,2)2ZJ2/H(J(TO#;g5(;(Cf
FC#<@g0/QIL\:+/AJD\IZgP&/B]#=5G^6+bEH;;A+:/XJA\JR2=;P>6I>3aBPVg3
DX[gZG#0C3KABKdE@#(bU@W,6L8?;&b[F#/V=)^;UY[(:WaG0U+3fE:,7KOB]g;]
\I[fF#TKXHPdf2&)V.@=eM5g-Ac1PaJ#9L6L:#=+&aaR05=;KAFYY0<3/AcWXVN?
d<PU-8Y:3UO[1FU?5(0G<6WXT>dV6X3)L#^G0M(F.9E(:W_a^GZ=JJRC][3R/1aW
7V4>5W[EZKUUIH>IO,O(8J[:VPEF4JV((,e^cB8.+32R42ePG[X@c7M_,X@^5=Td
S[9[QC:A?d_:)e9>@dI5?Nf&6P00c)91ZI6>C6de2AH#B@:J/<QU6ABgRM,Me1D@
^If.6b?+g6AOd?LTM7U.^0].X.RT\GH4OOF(25I#Lg^BYX)1\1B8?VC)N#UPe(3]
GSAM>TZAR;a<\UHa6AF4OQO4Ra)3]gXd0G6\6PGYXAW+D0c3,?3U]^A(PgfT=-]T
[3Q_P.E]F_@FY6MY3A[DJBQOL@0#J/6.-P:a&<+6Zc4LJ[+U/U?Vd]HVK6#FAVA4
JT:PCLe>SdSJ>JK/AJ_9dHRF&g-dZ]^\HM_H:^2WRc)N(O/\bL[4-3E+&;G2LfbN
1/LN1D6@+H4T4CJRIf@[W6P#fe0E&B>Q=8[U4e;._GQc,C=1:dDD6,3IF8WL)Q.O
eZYZGZJ;dCV7S6dK(-Z[gH^,gX/,G<0N5/(94I<)O/3,XJGX^B7GS+fdPRLUdU)V
JgIK=<J[XL<>1(f&KQ\J\)g5aCS433XZ8M<J;KG.;H[(H=KC_T+ad?00N,R[LR[0
0aaa+SSQ1IYW7EOG>[/BAOG)B8-647[X-QR;EO8Ba^E4;B>\c]C+YC68??;>b&(@
\8KLO6O<9(0.U[;=L/8M.fZ3d[.B:7650]94f2BCG(U,_GTAf=09K0@LcQT[)V-J
Z<ID.3.X#RXEJR\OZ0]2KM=:MaLd^a]_a;[<f#I[OHfa/P=>H(@<gC[b2#GN=/U\
GCV:UR08.=3U)CEVeWWGWR6JY5c,0?W0A,Ob<&^7EP3PYBFOL0(CW<67UGc.6P:1
Y?[JEeXM\YCXDb8U;gDcW[G6)N:&c_.3+e:#?K2c3/.V?eZMN7?(AM-8Ue]#B:LG
@S]QNKUKbN(0J6JKKH-^8D8=A29_(f2R-.=+&Q[B_0.X4SV].&Z#6&<+S@F5Z&][
J.5b<Z2.JU-/a&9f.6J=JH?Z\ASB(;AO3#3E+U_9WAbQfLB8@4b=Y;Z2D)Pf4,;Z
8+?=^c:WI=U9RBPaRL9H-PD\1XGZAPg+A9D@B#L0QEDV)OEN<VA3[]T2A.@XA0#0
gGBEGGRHG?UB]&.]MQe8Kg\,1K92.DEC[6gf_H=CXa[2EMCZKASHQS>Vc^+2\aV&
.2eZ\XMW?PEEC#[=_@a=/9GWd_7O?D6fJCMfVFH9;]:/I=6gHK7OXG54#eB.cF/E
H;TNPSL=&Zb:=I8]aSe9PQ@H<IgVO=:MD.^Sc;/:fTIO;dYHQ[/Xa71NJQ0TWY#9
e[d9?V2,-:C#PR#>cLD4@b@]<@F^Ff9aDPgZ-(-g9>fN_\E@)Naa/?WT1c)]+^<g
O[;Z78/4@bPRD\,-F16A>F>2e9_/YJS&d^&M_UR-^2)J3@F;_@\O6Yb6&6SVUf?/
7bZX9LRLW>L9;0)&,ZX?.@8>c#OAc_BF]Tb#gG,EJ]>L_JV3F4WNd0:L^K.2f+)L
\_]Jg^[:T07d;:1=a3EPOMJ+T-7Se&.2YC17<1gf[0U7627/)]>bg:[OC/(_bFTA
3fALcf52U\GKSKWe@F&/b<_WbO1<g)7WT.;28\g2TbJKaTL;:0;\4a]9=2+D9bV[
F=&Wb<]R/MABU4&STK)\2.4&I1_;X?e<J0f7ab(d2,J:Jc;S-A&DH8L?TVM<;.cB
d.PPUT6M0W)Q1JLe7PRT#?VR[T:[)]_S\YJ8)#[:Z5#f@16>LeA/RG_N^>Z]cL\g
T06DX5548SC?X[.<e?[H9+9DBbJVg[(ceTCJG-)LU[M2\aY^eL-@V45Y@SNd(JG?
;=+S8HcSNO/HEB84T/S>8Z5)XbELNa5_,.^1(MUfCf+^2=WJL6>AAf<[-.^IA@Y7
(J^).JBG8)PP.X0]G6E4Z<CEJ-)A/)fYa\@0KR4D=:O[BRD?5.fQD/>=5XMNVg5+
b0^68.)a(^\4_IS\6cHIUWEgc?YOAP4c.-DN<;-dbDZg&C3f6QaN9b)2CUP-Q:QD
RDg2^:XZS302g^D8-CZ@K#82TL5=,e;Z<_5,O,&&b8[J&aZ\>RGQ@4f+#E>c4S/O
O&5V^5>eJ-ZD_[fI51KN3.3^gOC?W]CL#PZXC+7T4>FRG7IK=3E0)(-N,-QKL/@#
2Z^NG[,)AU<Hf7B(:HgFHUMX:^e,YWJda7.]S9VR@<RZ)aKO<P/C2@.3b,N0@[\R
K5C=P55BY86YS8g[WW.F(8\@_H/GW[45<Pc,U)C\V+JB>gUOcQIFcNfYY_BTRJWX
T.WVB_M:ZZI)--SCG7:Sb2&-1Y>Fg1d<V&S-aO>E[V0agQF68L\TG32Z/S;gb:/L
EXF&51Lbb2.Oa<cKG&X6:)eXE<aD@7^S^JUTU3(MP<#XM[SWDRA^HED&R+=9b8fI
6&M^3<9F;R,WF^CDME38c#Rf)62#dB<E\L2>8N[CC]^;Ad&_U^D](V2IW9KT0>(M
IgVEBQ>^B104WP^O)=A)<Y<U#W&J317\;<UK@[)6,]LZ;6@dUCg[bQa];=NBIgK>
FG/DgQI,7Z1Y/O0CAe\E=&7^8=98.]Tf^g>1827[A?^)<dHB7L1.a<>3,K,X)[HI
3W^^>3I)-?R@)>E0c.eQ69[WfV-LV)=JE.VZ+5C]_K[2&DB-8-Y&N_FDT1JSU1H#
JA1>:-5#9I^Y]+J3PS:9G5,ANFS]2/PCH+K__MdHGB-@BTLNB4)#R.HE\5-Gb>d<
_S=2ZVR)1MYI@_A<ZU9Z>+?U]aWQPd?d:[P89B7e9PAV7CPAJ4[-HXVb>bb@g.#<
>K+:^:#CgcQ9E4.aA=/)b-U,B;:A[5c_6V+:51TCS9+KULKE0C@E-^&_F;cU/c]A
GGeOKNQ)cX<0[bgM,7>OC[N<b)b6ZDMgC:XSNgccK;LX.2^C<9?,+ddOG3<\YH?c
&IZ^XL96#^g,\a7>4U=&^\IS/IU:N+<aOC(YVK9?JE_c6e/(;-,eEa\)UZTZ]JQc
T8GR/VX<SD@:f(P=Ff1O&eDVEH?Qb&gHDUJ\0K+JI&M.8.QUF6L@5\?^))#b2g>-
TML8/Ue&--W2/UQHHH/TUWSUg;MP#6[;>>97XVVSVTLS0F@^.Qf?df<NT1KR#48:
\733NaUJ3Z6ZWM&Wb>3LKJM-@TMR;IR#U&^P)/Ob.]_GPC8@d39G0?72B?6TKPMA
@X/^)4R.7-e\DJX(Gd>X,Xb4Ha;f#-JJO-efdcP.&JYcaGXJ@G6dL(_3SZJR,A\/
P6U2)a+[FVRa_1-Y>.]ZO.249;Pe+)O0XC:[;(gbPHV(,OB#D#(V6=TXb6U(7d5N
H5=M>/70f<6TX[;WRI3f?Z&&VBg&UCRN8:e(2P]X>M>e\/;B,3OJ]\d?f[[86dSC
g\,.&3)]^dZ;_G)dV&?Ndg/9d6Ie[52;??\=I<R+I_cd8;&Yf>.<Pf,KTVb^-g3K
/<+0E)WBCB#@LXFS1E.P0,.L)@N?W.WT,d9&>[f7SJXF,=1FUJ_CL1])W?WGVUS>
,Of#IUNW.EObUDLE+_.LR)bgaVcQbL=a(NRPBUWL8DK/EV8QD56WSC?0[GKgOYXL
1L-QaO)eeU68N@W7?gI0VcfMGJPR0M94&0EeOI+0B(J2^\JNG38X4^GSMBBBK<8>
\F:dH:XN4DR(F,ZLW:^F^T(KO@=FQBg/R98<<C)EVgWc>G2CS;,Pf8#4:d=NVcMG
\1gG=0<Gb5c^QQ1>6FK^/IgGBc#(M1#gN4ag@&]b#O174C_H/\>2F>Xc#K,aXAT4
?e-JP@DVQQ0.)PJN/;7-GIQ1Y@;)Ob),K<.++_^GOM&(<3b/>ZS0f;<a(Lca5B>&
CU.@dL(@9HILIQ(D;#(/N#AfN+bg4IP7AA\fe.0].X+33)3:/8S+.9Cd[5cXI@cG
d^6>Z[]ceS0,@<ENQCB78(2?77=F5EH]E>MQIVCVDW;fF(EcggJO2Td5,T\?=N22
Fc;KMP.4fTg1)IHK+-6ePP)-Cdc\EHCaO=L:;\6[W4gbJe(Zc[);/Ve2G1d7VZL?
?M0g/:+#>T.=/D?AOdR<60aUZUET2SDD)0LQ?8Ib,0F\>:_HJX[,Z\+(]aM(K;cV
37a>dO-4Y2.6XefHJf1:8^8B]ebO_HHc7/-Q0T0T3TZ[BAKa_0g9,;DZ9Z/ZF^K3
[=C\d]Ia8\._B6CNfFe>N6J^.YICHWQ7-O,;?d4M/7^K^a):I=7VEXaFYe26.I./
Eb\V_FOeINY@(Wb_f=>YK/DLJ@/64RD?AM#=]DGEU<NXAS:gU\&2bDd?7FRd6+W8
4IOAA4[_Q?6_+?3R/U-_Ya@V5XP\&bSLP>;O+[#YI?7T#ANaJE0WBI[\9e?NUJ&5
:ggI]F&cR#+(B>fVD1D2)+#76TR1cPBX2#eD(b[B3,D4-34K[=XX/NU.]_cd\)HR
&+G)E2N+5#PG^=d470dWQ3\IaX(I5@X<4ESO[-CMZ(.@=@c,fW0]/Vd@SbcBBg-W
_-aFQe(RU6TJ+(KA9f:,?QS:J74KSFEIaeDF&1ae?fCZZ\)&^5S>N.]FdHH0P8.U
<XH8AXMO->N46LL;6TF+^MKM^&61ALgWDaD@#2gQ;_:2G_A5bBEY>0+]B)O)_AC2
B_;,#D2L]B2Kfe&\4,7e951gBQ_YZ+R4#]T)5XGC^JZ6,3)Q+J)7D3JW^T)d[8,a
\E4KJ)H<ZO:S)2EA>+WJOK^+WX9F,K;JNZ_1AW/HD@W&TO44e(X#-8KTB&;)JW8J
V6(QL.c[5EJ^B<KbZHcI)-NI,8H^.S[OGZNIJ1;dOXQW[f\E3&;WefP==LM62bX0
K/cU[,AMI1-S;O^bg:]d1(^gII/3,BQJb3#Egc,S^eI>Z-QfBG853TZYREMBgH9A
YV/AWRPKHS_fF2gGG758FVL[Z_EQ<^(8NLYTIV#N3aHag6+PNNg?gJK&g3DR5)UV
L^70UJR1Tf,CRA(#&U)\fY/ZICf_T+8WYOD)2^-PX9RcJ9Nb]E:e:fgb6<NXeO&)
E>,DYX6RK&a&80\_#AM@+S:-FY^1M&_E(YZ82B=AB[JYX&LQFN?(E+JT9cVRZX)U
H3)H^6AJ??)0g-BRb3<8_(Rd&1SU<eX<b;>)ED2YHC7UR#]#G?,)=DAMEGR__-gM
FVW8B.EIfWW332QPOPUN&6U2;&&f^dT?3&ME.1:7b>,=Q<ef]0f4#77=K&f\>(77
AO^L7F2GS<#8V6>HG#XTV#g47/dX92-KRY?21Q.)bT_AD^]SVd@&6UB:7<=I(ZV-
V+^R029:,ELE&fe_M/bP?6?G\#)4#)3d?<2bNgCZ?>9S7#a0>>Q1_^P&SJP.C18)
?0N]D&0+c^0c8K-PQ+AE-0Tc>@E@6+Ie\>K>OJ=<#IOEL,SAG4Z5Q:3O/Y8+d>>f
H/PM+fA2XL#W7XFVb-27e?J6FSM7<WM9N;23J&L.JO.;QdE]CP#g^I6E@&[R)ITT
fHK+bS@2A.)>aY+bT^cEW1Y3_?dT-F#T8<+X[V]:]&T2Q6S/:BBP-+(N&\#MYeDI
3&R(-f-?=CIc?7JP1,L_P;FV,#W;@JJ;>&@P[&_T,MgWSI-/)=G^Hc_Q#ET[,4A2
DTA./[c/B0K6]U=1QSJUGAK)Z:57e^,X:8Y&WX;(X]Fa_JSSXVTfZ9E)9+<T4_I5
XI8:Q^I5_FHLO/H.50(&N>WC\B7F(A-[UOME&#&gXd9EXIWd0??TW^MSYcc2E_7V
67(=PgF,TZEFE[eeH5_EGN::#SJC4[WM#Z@(8WJe,_^Z^g>T>MV-eS>C5_7fWM6U
R_)0T=XWWOGdW66[SgSGSe24g4=WBdP0Y]-;_T=W+&eE]61;<_N=R)K?1;b^ITP7
TF1D?J+(fXOP?C=CF@8)LXf&bgaXg&M7H_6YAQKbH_9Z^<W49YaAIQ\NeH(Z8)2@
\:1NSgCMN=S[VYPP_/7^.]8/=.BQ]Fg.f>GY_>GNL_UROf3<IWQ^Q]YE6Ag8Oa(B
de?QK#c-7K4\HU1L5Z>9]OeP^41B74a1\KH?WTe\H^2YOSOWJ#\)c]<1db5eDOfS
:7.F&;BIMN;_#54gWR-=D^?Y_O/@&gWB\6#L)G8X=L:,YE.(L0?;.5Y/7I#QdWY=
H1MgV>@GWAcdTKe[\BgcYa_C-;/#4X)QIa6bEYcJXS)Vc]L-;Z1b5/H?_H]=:e8O
5R[E^JeMT)#e])?C;>Sd?-(_5M\dQ@I0.>VRHGN=Z?,=V6B[Z5:[#g11VN\OE70<
-OJB>9I>J;c_/86A27[eg:@UaecSg/d[A(Sd9>c7GWGe+4LG\B?>=3GCHXfYVHBe
MJ3aNeI^bM20TQK?N(1NBWPCfPZ];F8:<C<6O-A4[g^ggdOf3NLK+&(VD^D].dC@
LO8f8SW;eOLV/fIbS&Ve&;/];HZ]#?>.&RT\.W0@1-eN2;)e1]f(b&+6IfOQ^gGC
V5_8?0:2efD>^>DA>S^/DGLQD:XeRb-gBF:Aec2)C>:#<^JO(b[>[:gP];]/#3(9
C?bJ\H^ba2U,/C]GC)XTFaJ8_ZeMSZ-QBO4eLbGYg#<Wg[-(+/9/L).AV48;J2Zf
8#2@56?#5[\II4MHQDNRcV:H#V_ADHc(,Kb;.X+_M8Kd[6&gOK)MZbcVU)SHdSGH
@7>bH+F./dM,M)H6egSeR>1Z4Dg)/Z45cO.AGJ^FAICEWZN]_6\)]T,N.]U:U)8=
H&.2EO3BPa#0VM9B8./X8<@gQ(\5dbLcWPE--AT1N-cP(F:RAg(1cDU_d@,fV=A.
M@+N^#deAZ)02Q5fS\6g9#<We-&TX+e^H=ZYQ:GJ4^fD@5?A6&O(;f.LCK.=F,)2
^d7HD<M\ce[[PC9]G\X>?Lf?#Ad((.YCg/#Dc5#>@;IeF[/0Z(HbbBL2_<,DDQ.L
R<B4/EPP2F?F1M+7ZJG9<=2.gT]@Se\LO1<:8AIEEDII9+-+(PTG;G8g,/Q7W+cc
/I?Rfa-82GKY,VB1T2-\R\4DL;T\a/ZA\_;^+PKJJ#J->Q(b_VJI+Jb]>3/cZEJ?
PC7U0B&@A/G_^16fI61#4)4#Y1Lb@VNW?SVORVd2JML=ZJDb+6aQ,T#&W3I[Q/cT
@#F^Lb[K.M5@R<GL39X]BA@08.Z\RN,<1KMR)+SDffITH=;Y)3]_W/[Z2K(8E@Z3
&cK/RT1XD]<\BRX,E&:8QABAb5QZ+VY,7)8_ZcCdAPB[f/WDVFN\]5e>4a.93ZeT
YM_J]4[[\\(R>aQWPf[NH:>\X_^bQRHXNb2e<SPDC6MXL-\JTWD3L,g\=eGNIda]
&&4DV:/GJ_MOF-,9D82ZFcdR:I7?7^g253@2F#QT2CCU5Y8FZ</GR<8WDb,(?Y=?
cQ6\\-M&2J8U?a<]>5Cc+O^W-X5K+@.;NYbB(6V<9\d8g@AGgQH3JN@5&/:->U/8
/0Q]><S&WXIIdWW<4INTGW9EGF1W8OQ22]LPJDBU=5BcaCfV+\C]US9=AFO^ZZ@b
.[@V4R0Cd-0UO0&f,^22dO+4GRWVR(0c15L9<,b4IA&9>\-PT_:Y.F4:2L]T:/BH
7R;&4JT4@QX,MCGNNI[BOK6T5^9d8DYI-e6+O@HPeX\PB053S?#XZ+YJ,b6e.b\U
Q^CCTR-[1B<#L4:6WW\3]d:WBf]AcJ+:H\8gXAV[DU?bK=E)^cfJ87(=RJVc=T15
=1^A(/R,SeL#@RJ/&6Q4RMJMD2BXd+R\.TUP/500[N(R+HKb3\cb#d30UZc.-CZ4
4T59^Yb++&C?[W4fG1CXKW.(7HC+/XP+/,>CZfO^Nc;U[C/:.63?_#2::EQL24NJ
1GIUW\GY>(^9&DEV:S10[SGQGe<4HF[9#SBJ+FP;d29OWIe93#RH.2dP<[?)YI_,
<[Ha#IUKeA_Z@_<2de:)O0R(U;H-8TAR80W>O^^DHd@Xe#d)\+7PUH[8X]UVO,+Q
C-;)PD9+9JQB#Mae0Y=-/;9D]5(W#(]@8WP-QgUH[T+4SW]5a.7bW)@C,G670]_[
OaYG23(?(.)O.9#NN>#+V9I/2,Ic\=YTDK@&AR7GdBR0D:gf]A)Bdc,aJ#aR=L0S
_0+T#UPd.)d#.D]A-RI+TO2>g\a.;I?HMN;N3EP@PU,#YV?L?^+3Qc;/X/+a>dSg
1IeW^I0(#9T6_LXa&&V/1Vd:G.C_A;&J)7V.K[Na8[#U(DB1<5P&.>C_:3M1O6<P
ZHd>0dB.+RX]\A8N^,->2(Gf@RDFc5HC1IQ_(W7VA3egN_5(SS4\U.;?eDM,e\YT
a=W(3:OT4+CV)S:38P<#K8YbKd[FfV0/ZI(e^RQ<#M.BU(T9-.YG/F58Q4K66A1D
b>O8VEST:e7=;VWgE_=&[Y1-g32\;<E;QEVHM\HB#0e[SSfP<2[aH[)MZae,0CS3
b9T7A+=DQdBBQIP75_9Eb;<>4CRb+GA3[KX);b)APR4(9=Q9_JVRb=V:[)^+0VEO
DV[5(59/9&Xg]X6;:AJ9)f6IG/I74D=ZYAZCMEEYWK#Q&-2\f(>I:e=Ueb<@LeGe
B>(/^eL(,QE.Q:.&7;aS\8MX9]7D1K#S13___)>1_=L-gb7H5GLKW]c:E;23R9T5
-Ye8,FHQ+KZ2O2K[Hdfcd>P7Mc2?N3Qf94K(3/[147#+TEGM8K(,.6eO7=aCcG&?
B8H1_D<FBMN^J?;9_9435>a48VT<M516-cS\f,G=gc</F/@3H]B(/(_IU@Q>HgYQ
C(f6KXP<?T9/,e1bGEf7KCYW:(b:^+R;5?/DX9?>24=:V^Z2UHDJ=32C0C3OQGX_
d)KFVc8A^L0:6T=bM<(KI&F#PV&V,R5,+,gEb^eB04U]44R<ME1#MF<AJK4c<0AA
/=bC)IgdDPaN,B;X=,WUS4/[L9LU+/]EQ2BK^J)Ga.=gDa)\FY86SQZ\H442GT(Z
>AA#=A:4/ZK2ebSa/FC_S,fP:U+SHA>B;aJWF36M=GaTIcB[D>)@^Hf>[YKO#BH,
_NRE)ac+W&eWVU1f5a=CfD<.F/KbV2Z=V8Z>JW?/N#(37JW_.FQ(fP[(2+9aMNUP
ROCHIJFO/Wb+JPC367\H;O:HM-4B3K7-@NcYdFYbZ<J60\IDDAGI@DBfR+OA,a96
ZE>&&7E(dYUPEIDR);1XVE-L_BU[eA@<=0?M[>N@/f;?NaP^T3(_ZDOWL9D=^E^,
O3N.?FVe26OMVTT]aP7Wg1L&R;W=E7(#/2@[^S[7+F@X841NU?.JeO[13F]fgbAE
,&[&:3PX@G36XEVae1^V&J.0:=\814UT?2ZM7>H)e8I6PfEKJA,TJPO]C)_NU]K#
H?Vc&_F/D-&M2gM,:YQ?Y/=D6HN8AUJO[1GT)fG8^e3OS+g;]CPZ<[Y8;N8:eAeP
PQGRYaN<U9,2]f7YG\gEPAF^3+J\fH]2D&NI#,3DbReR3]]C3RZ5OVH@=1&_RGB0
,YAQQ5_R/6:\-/-_E.)^.+JCJT=PKR-O-X0;<c?\Lb?#33(KN0XKRQ4e=0La62L?
BG;1FA@4f;aHG]/R2f,^G825GAIT@7b17dD[D4DJOb/[>(Y-(D#&<Ne]dQL#D2Og
SdPC3W/QdUEJ(OaIZ<^M&1e)O+^,L\0FW3GeRE;<?EC^S#8C[IFb8eZ3J3=aDg9e
N2+;F5BTY&;[BQDHL7I;#Z[e)c7>MNVOB426g&1/Ae_]9Rf#6E,3fA+=EId54#@O
dQT[U(?7@9,=dBeBS[L;FYQ&QI&EU,\A(ON?Y3W_-V6BL#bBR>(;25Y;[F2[a]+E
2TB]MB6gGD^DD(b6Z4<S5VFe_<(1JJWUbPFNGYN<a=A^6gJ(N;8faHNeF;(GVL48
1W8LZ&d/=>Jg1FLQOgWKV5C.DYJJ9\SIc4:Ie5T4#5_ZCF;Z8=QdGSMHOFL&@TY>
K1_=#;\GRGI8W#G2>dO=GLQ@AcSV3b33IW9D4a3]REP(8SM=bdd<3Rbg.(OS2CgZ
72\7_9\7C-(,4P\+LZU[ZPfN]F+@JT9+<#:,F^2G]d5MT430VFf(f:2K5+GPg6bC
CRV^USJ6L=D3aIC6FN.Q=6X.&7ZCbCE0CM3LR4WBO6a==6^[RADI1CdYWG;=JfLK
5)16C5@1/<[a)Y5Q7@].KU)^ZS@;#gNQUK@ULW;1TZIA#.?9R?]KC=9C)&AK>NQ4
eb#f-N/f@8(XH6Wb@0?(W;VBX\/K(--9_YN/I1R^.NDYTH7:8D)-N0>9MEVX>[eX
f5O&WJ:_;^M:U10Ce0C3<ZcXB2R2OX&GG?9Q?fT^c/;R<GWe.fNgKHdKQ@].G59H
NL_d\,d;45_<M)5R@JeK2g7ESZRV(W>3;&7\;7S6JebASF[YNMPe&D\K.3HE3T7_
6HVa5G\U,;f?4,5?d;?7S(9bDfC]GQVLQ)+2-Z:?.@Ba50@+a;<SETXJ,Z\f]DC6
[FX/4N6<>LU:aLO;4U7(SGZM[&g01bDQd;==aG+2@dQ,L^,I4?d-])WVZ:Xa<&#B
+OK,+U4eD5EOSU558gVQU^@\N<+L]b=16[8DS[G<8)/?S17E#e2Y0KedZ?-4e.=I
<Y05bagYB99KV0ddf=fMU+WE:N6P^LX;#V+L=J=R1E+QLO1/\N,-cH0LgUf(cO+1
03R5982?C0B<Q2]XR@OO,9,O9+,Yd&&:fN8>S.WD^Y>F+C0?]^@3&@7.6B<80/?/
f380Q;Z]((a8M>;)/7VX+13N-N0L>E+4]Ja9/>+\(.<J/QIP[8<O<77+g]1/K.GF
T@^1TB+feEU.SC>TWZ)C4=PJT4AMK=C)f:DO9C99B>d6I=]=O8Ib+5<M@Z873CAP
GL-_V-3c3&OWR2J]/\L^MS)]+A]BTKeX><OJ,:>d:..A4Z2(HP4b2WTfK?@bcJ=b
QDff#gG0=B&YN;(IQfI1/C0[NMR.&)QaI91=C,ISB46:a2\D<?K]B&+9GGF-QDIX
^dU4gS#I<)3JC0XSGe_W?)Sgc,gFQW3I1#E:d4g?1V=NK>&N;_Lg@/-QIGAD5(#g
=aM5L&GZ+X=J[3E+<HfC<KfC-Xg<d3e7G9-R5RO#/>=L((EA(4bc+KS>@7bSC8QK
5X]2_NM+M;e#C<QHI8:8ab3THTAA)e_5S][b4\NJM3:;2g7b=HYLNR:,G#eXX=V<
eKB0?bPH>,;EV4.#.e4)eJIcNP4I=YcBJ>WRO0HPe(:DFV)+356W881XC00YB>@-
BAKU2=WPL#1UW1L>aec&@ge\\A<_@&9U@((5QM3ZXHNV<6\:?a8+81OAaZ;WeOFO
f;SVI/)GLeX],5E=B>X-1EF(2G:UWF=H4<4PZ;>XAHPW8AX7Y+OJK2.&U7Hd0,A^
#:K&=>.JGf-H@0:3^d#3U,8PJETNBdYM/K@^E8(]0DVe7c?^A6IgM><4J^dW&H/2
7/)8ID;;WL5#51L6=KO_(YWN6g(0>T+_1I\JG+_),JHWZK&)YA1M8IG;?G3_CSZg
V,28)ODCJTHabQ\)M==\+K/^]/:JI(T>=J6L,:9P^IQb3cY.1eS.I,,C7B.ZOZA0
11:5F;g58]SB,(/bK(@SeNUD^C7[d_S+55Z\:N\CS9&.)17^M8&2BF]VP2BS+7)c
Pa[4/(=@/W/Z=f+J3O;00<eBd>,XJ@5HHMSf)aaf^,ZQ:&JD8NgO&,ge97edWJEV
88D/81O3N.M?T]c]ANNO.d_2Y0)Bbe)RRMSECJB(8@A1XY\FF@N+XQVHXbQLCC:f
8MLc2(6F_+##)Mga84.&@0=O-DN7ZUM1TJ8CVV@0ge1+OK3G>&>T8M@K1JLY=[CB
7>&^9e6C4N&JZ>8+OTH2bPaHKD7aM7ga<K>-\6O^#3481[NMT=-AD-+)#C15-DQ;
K_D1ZS,BMDR6D42I-P=H,b(1C05Q>b=(4KL@70[cP9(KaXH5(Qb+HA5EN;AI)dTA
b\/fYa/Z=GC5\A2MX9QCd542VFU.[9[RgR&ANR-a^Y;e.(=31@e=L?Id5Wa.B>A\
P+?Y,2fAD29T0d,2X-J)?#?6SXGB4PVUae[O2+6RgZ#7cH<OF=8TH0USW?DUD.Ea
U+:dS[(N009,]F,ZfPb586P&MC,1@_:_/VK2UTZK9KX7,c)IdI9dP1<ASV3fQ)d&
Q:@#(/^K8Sf^X.bX]LA3Jf7?6L_VNLFLIBM=C2K\+R2DAd7;e9,GN\KRd5Y&<S;:
#:?>d]DD237\0<H6-)Q^82P9^&gJSRf4?7LP#MRP-583]FgW+@T/g1?6gV.C+?H2
gDCTb_WbU#FaK)Z54?>.Wb\=&4QWFc_D[LD@&[]/JO88-\D;I5[.2edc1QL+/d_b
U7&R)&R]GZ_b>]]PRB8_IadLO3>D:+;J8J#ZC.9M>cQ?N-PDf92We\LJM737Vf]7
PAL2Ia5M5fV4&6Xa5#>WULdg1M/C#,#+XKd^\+1(c_Jd>;(5/&GH7:ZG<^O-eD?Q
M3S31XC:Dg;a@?8]U@a\/?[:FQc^Y-eIcYSKU5O61=6I97>PF)b8UZ6L:d:3-0;W
^gB^6dDB,+[J]?A.91A?@P+1,U=I?=5Gg(JI+=/5OVF.d1<bUa^12;5#35KIC_+D
4VKTMg9K-H0A3e]PNZfI8dM01D#E&1PX#3dUCW0LO7LCE8^:8C[[gT](:F^=5_(Q
18NCWZf.F3:D6?I/CS.]]P]NCa+b._G)S#D=,0@A9.G5#g,6_U+&.AT-c.Nd9,f=
5BE[MC).VK=,8KUg.[G68;XOB5_H]?.MKD:8/RY0e+dIV;9ZYa0YNKbU@f56K@KJ
Zd-9A+S0:#f4)/9_M)FT]TB]U]@aJ9[HW=?KE.I:GM\HFdD2@&T&/+G<Tf\F13Q(
L.=TR1D@KU+G]Y&T#RH:?-&;9UY18N[6C[+2:)/90CJ+cTg2HL]VEQ8.Da2U4e[L
LFP5ECH+.-3Kb?S>d#0U,-YY,ED4&<9-)::M>SAcB@_f:Z/dc+5C)ZbDGd>)Y[fe
W4E/QO3e43Y31ZZ&@_WaB5N49G,B6NaV)N3eF.-IUg5b5;;Vf0@#TZFfF7VW8b+B
2[:dWB?=a8DT7JDSIP-HX:,d:85\H/cc<aJAZK;A(:@AV5B&1_8NY\[[TcUHG4BA
9YE:eT:ec3#0-bW)]E53X)2_L(N8XWG()T;]@OY:(N,@5UPVWIf]5&7M8-+D0.?0
5FZ(WI;V53Z&A&V(=M;^K:beb0&f7T+U5M<cJ=.M>?ec\D@fXJDKc,>Pb>dGLa([
JN7Q&B:.<Vaa?<F-&9>1#TWBIA(H76:L(JgNZHDJRX0?MAY#96f/0PSSfEaQFFC\
@#R1:.[3TaEMIOV)IPKH-8I;/;g7+;/2=gB=GF#bb7H]>bX4>?(f)-:QFSTFZIPK
:Lc4+Z>:];>SF[SU)Cc))\:&KFQJAOYZeZ8O/^4U8Zb](O^J^8\3Zeg5<)1/d^^a
/;B(4-FZ=7SgeI&,>?9L:Q\;<IS3T.Og#/0CNM8E5MU&D_1\+7c:gZbUWJf4,W=C
BK,#C<4+7+2ET8I2.XE32,ZN\2W/\=0IJEEP7K&7;F2-J=\^KK,RVXOg28=786Oe
2UL<D=a[+M;/OSWgF:e7G,d2=:8R<G?;OY9E=.U:b\2aL+.[C7Y/R/H<K<E.A5E.
^c,:S>fY#B)EaNMNKCAAA5FZ#g6e-T4P#H5W#6fM7FbGP;(_.)@Q_dV9[EA.P:f9
1]1SY<;UEX5MdUM1</SBQaD3?^@,CKa[?VUdd&Cb-ISWC3PC4C:9^4Y:))H/cCcO
Q7T\:T3b@@(GI_OR&-.\9JZU-UcV5#RON:6&:O#T:681cKZN[XA-+_L_+IRF0PF)
KATAX=BZJ.WW)9D5ZJQ2J#cT.e1R&QTFSfd;6@-L>D8gNe(F:@QgT8@<M[M9T>N&
L;48O[H_8[_5P.16U;L@M.^?(T(J[fAR<e^XR]3(ScR[FY]RLC9.DMZTMJCQ^.+8
(24fQ[@J6ab/14SdHT:N8^1Q4DJQ@+;BT.IeWCV>X7R5A9aP4J6Q](QX9fP+LCZg
2<VN^GP@Y4IA;LHMM\c1QUQX\_J+#,^cM+G2[Ff]IdOH:BfRUG00+]XE6[](RZYC
c=Z/15_D@C,3B_TI3Ac]U<805,,PZc9+->O(>Z@QW9/d_;#FVYMPaSA=1.ZEcQ.O
3DEM2DX^Wb4V[LgV6G>V/?0/_?Q?3E]I3<Q+17c6SN8ZKV=K17gbgG1>^9IcW=RM
Hagc:PAWI3(BRW7AU/?RgDeXW)19B+V(=6Ec-]X#OB9][cdT<fHOUYA)U+:]8>IF
#.\>H)^<\+V\QWU;6Z.8P?#0[>e2d[6f/>e@701gVQWCH<_-]3I(-IGT&Qd(=VQ]
]Be>.fI-O:D++]g#5Sa5WQYG.8&>+Fd:]U-8BPM/+X<[3)H]=7c,(Ea[@E(H]^80
JVCIZ@:IF)[&FJ7E5g_@1FJ910X52C.&8O7#7+0+-H\R&X4_;38Z_#X)6W#J\]]R
2PVcHR-E4DUPFVR,R_QVgKaXD&=)51_2?CC@a3.D+QGTK),-V2P9ZX82UXDV9NRV
26OE[DJY]<<eM5O.7#Qdcd1IUB^MQLHS_1cPCTTa:86TIU(7f5[[3B5@OF?U/[X9
/gX14=H[cO0gGb&N-CgVE_QWS=ML&L],K<Z72@^9-+DX8WAAF7[#2IM@@e^(8)BQ
a84T.+,gZ5>>_fg^9=.I4VGBe\LZ8IPD<6EeW^\DF5./-8K+2M)YXD;0<5]3K;0W
d0^M8O@?U_=2>+&;Z4eab>+L_DBf-a8D)+PAU[DLCV=_-/#]FN,SBE1\-SV\]KRH
g8b-ONH+H.8-.=:.77X:RN^3Jd\78>EBIP:#:AVF#553^DY?9GfH;K1g/-/TC?R5
OWSf@R<BX(@.:=A>G(@#7.]+6N9;C>QLVee,MF(:J]>XN@^BRc.K?UZ?SYNK06LT
F,af@^R]=f]aLY(+1^72GR1(.&7:+U\X&fY3(AN]#:<RKaOR=0d;G+#@2/gO^2b2
SI7=30#;Ef[-T;OX/</Y+JW80D=#^+2.&DgeAQO]F=X#WV,19R;HM?QQLF>O#2UJ
.F<6I8>(#c_g[I5B)?)Ke];_52_FbR3_4>=372,V\=-[gV1GN))_UO3]M4#>gDRL
-EfVU_26V^2#[D3&;B(P;S]OdMf^2?PL?#f4ZKTRH>;.TA?>L(=D@4/@>;.WTeVc
0)f)HA\0MO[9-NYdIdQGHKEH\Vd,BY-P6eFOVFL9.,R[&8APZK029PV4NVGW9K6L
2ebJVK+2Q?LLdN@d>I_TR+><-H&Qc[;FK_\QaDEX6S-@DNN<XJU<Q2<\2RJf4^O4
-<2EVe8GMdLE?<;g,7ZK2Z\J]&EGS/UVOPbOD7[V:3C<Y_]R\a]aU0<JZ19e:A3.
595_CgG7APWP#A7#Q-27R/3g1,gI1@TOAb5:2.-,,gHOda5X5TBT8];U_FP0Gd]c
L;)R-0d#f&:/H10/QXV>Y:DES._QB_gd@R2Zf:0dJ_SWdJ@N;.\1R-A@[JEfMVIa
#Ma60=YdES-<cb&dK5><V40e+=d#OD;@0(#:@_#bJHHAD=eEf.0BVcae8;NLSF73
e652<UbEd2A2O9F]AHUZ;,Zf<A?<WO+Z4N8]e=HKZ1RAT/BIYBUO7D8D+G\]N;98
bd+X=38NZ8g;<60:2X^QC[eN-VXcJJ0=-UVQBb;>VS#E.fb5IWGACCA,ST].g?WO
60[8#-dW6I6;U;=&XbV2C^S-VaBZ/\T)LG?C/2:K+>9H47YfOLK0Ze1?(eZV=_5\
[?)/+U>@+T&>GCFZL5b[bdK#UDR<I1@WJ5S[C6B-A02&22Q+eG#?K67[B?W9.X8K
-I7J@.?ON?+5++\^,(.-W9V)_QUJ_fU-6a/S9&B0LNbWfW^C_MB<,U&:WM7D--6Q
P3CKfRCU)L=_K-XdQQ#gd-gg1C_7<\@)NXPa5G,WGI)13MEad)e2DCB(?gXEAX6R
:4_N)805KJ)cJFD#Y7dc^X^SK)YMI/d1de?a9O8)@_0NV&1)#<X6H7F;R#(68ff9
GA#ZYA0ZKEXBA(LCA_S98a/51-4)@3bLK9OWFX[fFS3;E(gW7D\]WU8BH.N3&-2N
+4ScR=@+Z9#4]QF+c;G9R?T7-\,0+)-J<]4Q4eH8?D3gH8f#HYe86[O,#Pbf-\\g
.DVR4<HH-0[^/Z(WeZ]8\>]:TGNAF3Y]:=gDHXWY.3.D1CP]IRa,@O=-Og#,@HP7
<Z\[:_OPe_,;ZTfEe38(Y@F)?Z2)J->@a&2CYf]RQ+4309FD9(E\,E[08FXSLXU9
CZXNLRCaJ<.dH/^aX#dIc^@L/8(X_-6eNX5c?FC&,TFZ:dC1QGGdGP[>8K\4,T68
MR\ZIag;2R48).d\UV&f#e9UO7Y-^P#-^:80,<9_5((C+)G?MG9V:M_T4&2@C.:F
=C\N-F&0MFGI#D5BL1E.aL&;:V?9ADgd4O\>;;:4dQ_RL,U#?afaRT4531TPQ8VE
1VKbD&3Ag:Z.P82ZJ<J&^CDDS/0XeE)EgPHK0Seg0,N>6?@JcbLF,fN^g-(3HU2&
E264A.<c3fA\QFC5:?KG>G6N5^/3-4Z_UF&045[:PZ&H48,bU_BLHE;aC_\V6?N-
G6Q)X7CS#;8#DPI))(2ZFI)^Q>[:<P.&.1E^#]N18MT7BL.T-Sc+7aX#QXe6N>32
A0<-M05+96[>(Q@_S&_#YA^E,L)Fg1HUDUB1_4)7_BHd].[X[V;33c:<G.+JH#\R
N_=..[gPH3]8NdHDf7),OIU#AbG,1O(J.P3R+4A=IZ[BO35T>dKg@95Y3:NS&<0_
NC5eMQN[GU\,7&2R19,/5KZ9A/;EQ5]gE](aR5KOPJX:Za5,:]GO^(B<]e]L+G_R
DH:-#eI:g7]-)4A(FRNI:?\4Q]bT^&V#\46:W_BL^\-MfAWL7I2UHHgXegg&gcI\
OeO3Hd<FZ^)>-ebbP_aV,)\E#AV4S3QC[61\5fc8,KB7FA50/,W/[c[ee?[GE_=X
[D__dRW<^B@R#PBM>KYY+O::1UI+KM:(.de9<Ge?81(b&2E]0?J:6->DT72HUe:f
S73CO+?OAdd4WCS<R<Y0;SeIB1gR/7c<b(;](KL=2.cC-F=?)(\8TGJ=B@^e\19=
aBCA=a2C/,ST^O]14GDHRd@)+(T8VbC868,OOc?F&8GQ=U[CPXP7D;[Q4U<+5I]\
=^M7-I@fcXF2Bc;DV4(a8[cOA^Q]@?4^&.3aLBbZ<Gf+#-f/.d1dMP9e>?S9?=MP
QZV;e5<7>cBMWCRWC7:BgYD2&O?()cA0@<;CcI5+TZ@bN2&\acdP?,HDe7NDeY=P
UOa\P+/<g.HI<S:((LNJCb_WF?@1M2>TaU_a:C+=)VG@K=d:)L/8_D,/I+Y>eEb=
WSeQ1>Z@NDTWd=Y2?;>g7:-)d<f[[-aXg=15TJ;QR>&3G+LN-NKAAK=AbAR3)P=)
=GaSXRT[DC-9=:#>J>NR1:],5[YMWc0>ZR^KTKV=eV2GNZfNYR.:.f3DE[?DBQ_#
>HCR)Ub66G=KN3U3^Pe)MEM@:4PU0(I4[aRV.=a<KQab_=Q8_(T_+QOSYBCW9_R9
D(c1/SL,1T1<I-+Y20H6@?<R49V[f/G,+8J[V8gaO_\XM5;N23:DGDa#UcCZ&c]E
Ke?FV0\Lg105-IcRC8]5#ZNY&FaZ-=;@-;eZ-V=M7]J49_#WTIXHE+,fP?0IZbNY
CcT-((JIMG7Gg-#5&g/7NE/65EXH@X3M^R;Y_E;9ZXAKBV(,YeaC>J,&D-ee>4L<
H=>+5g]1TB)bgO2W6KQG3A;BZPXC].:@V>15_6]U?aF2:JGWG8(#6,eB?QE3-GA<
1cAZ#G<0HAP?9?,T11R\T(F>#FEc0S_?^1TX>#B2Y,dIQNOR_65F,93d]M<+;acE
XX3IZb\5d:4Z(eWP#[S.&J;,/d05(<[CUBK:>79?LG?7AaY,OMT+4CT5TP0CM5+.
g30R6/YR1;U8a9D>L/H/[M1+F25HP=UE(X9]<ZHH,<1A5Sfb];4/-<.^=/_[[?dQ
BaFX9DDXH^(4(1dHfB5;ZFg=f+1dQ+7^\UNd6AT4b5(58,bbaEdgLIW,X3K8UTXQ
;(_@#B6;dWVGg&V>:MKCb#L:[XXb+F</>UVN@<#+)4N1V<V1DE3@?P9@0KZeV;F>
[/+ZcX;UV3DTTed<e<DPL]^0VQ_(87WK6,E,[>e=12@dDZ[542<Ba,58B<+:Q7.9
(a>Vb.B#^T37cD;XXB?S:>+O=K;6cOR+Z#aLF]8GQa1&=c.F/a[3RRBR(>9X4JYF
]0bVJe9F7IR;+-gP=Q2(2I2NNf3IX06b4+;&[@_FO=gMf)3.f(W7RIfBOH\N&)T1
bS4U4NYf:=P3aP3Q:#+EJNV#2(X5@SS0IWLe,045Bb(,c5,9eONd^V1<T(#=+)aV
NGX.^2B-&TW<GM4C0JR9&cgMNUE-G4R)]VLdYQ,H(ZKab,#^0?>>bDbeG?R(T[[?
42.O7]+6I.D_Vd1fF\[fCS]e(;^aEUP4..=b4=EHWfBWHKR:IU]8e8[9E,29IY:_
S\V/f;;(Q[G(:8ZQ_fNCO:PgO1A^DWW4IK@@bG]VG,J6_4X\#Ja3H[E3XN#ZeZZb
0V<,6eO+G#C8;PP[WgXJ^=4<WH2F1AGc#YBPVK[<395@7M.RDTf\(JaHR#69H=T2
VLMIeGebZ_d;0ZX/W]Lc;0WH=Te=JbT(0>1NA;]6@P<f^)/d(2,^ffOE6G/K9U1A
;_26_6_e7gX.I^C4T;I@PXf,O)H3NA?OY)1PfD2?AaA#YJ9\>9cP_.&PI[(:_BIX
5-;fUY>[PZ<T)CVF#SS1E:bESgI-VL-Z\(1\fO67Rd&D5_Z];]S)UYSQ(PP)A9@&
?OFeCPZDgbM=,Y+cSdC5[F3+7/#ea3+M8T>^)+DLVQ0(e0>K-J-,R-]9F/f&2MA7
SC&;,7:5a>(@b.GA)Q>e&H>d[P?:MeJgJd(P]R0Dd_LZF4/NJC9HGdD8Tb+^=WZB
G8-M:_R/:cKP,WHN=ZbP>V3K>^85EaM-3F:2R^5NTK.#1;#D\B7CQIa7U#7<f9O,
QO8M:<fe_M1.ZcS2F3UaAQJSWTbFAK]<YJ1fgZQDaH^;&T1:F<fWe(DG<.:I24LO
;UMAc<R/HBG)A2Jbf?]MG]PUB;(3:\CcT)gFALY>ACgHgc8Q6S@&S<4KCAZFC)8+
S;g,2>@\A/?3C-.EAb,-GLPU4$
`endprotected
endmodule


