
VERSION 5.5 ;

MACRO BONDPADD_m
    CLASS BLOCK ;
    FOREIGN BONDPADD_m 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 62.620 BY 56.920 ;
    SYMMETRY X Y ;
    OBS
        LAYER metal4 ;
        RECT  1.310 0.000 61.310 13.500 ;
        RECT  1.310 16.500 61.310 30.500 ;
        RECT  1.310 0.000 13.810 47.000 ;
        RECT  16.810 0.000 29.810 47.000 ;
        RECT  32.810 0.000 45.810 47.000 ;
        RECT  48.810 0.000 61.310 47.000 ;
        RECT  1.310 33.500 61.310 47.000 ;
        RECT  18.000 0.000 29.000 56.920 ;
        RECT  33.620 0.000 44.620 56.920 ;
        RECT  18.000 50.000 44.620 56.920 ;
        LAYER metal5 ;
        RECT  1.310 0.000 61.310 13.500 ;
        RECT  1.310 16.500 61.310 30.500 ;
        RECT  1.310 0.000 13.810 47.000 ;
        RECT  16.810 0.000 29.810 47.000 ;
        RECT  32.810 0.000 45.810 47.000 ;
        RECT  48.810 0.000 61.310 47.000 ;
        RECT  1.310 33.500 61.310 47.000 ;
        RECT  18.000 0.000 29.000 56.920 ;
        RECT  33.620 0.000 44.620 56.920 ;
        RECT  18.000 50.000 44.620 56.920 ;
        LAYER metal6 ;
        RECT  1.310 0.000 61.310 47.000 ;
        RECT  18.000 0.000 29.000 56.920 ;
        RECT  33.620 0.000 44.620 56.920 ;
        RECT  18.000 50.000 44.620 56.920 ;
    END
END BONDPADD_m

MACRO BONDPADCNU_m
    CLASS BLOCK ;
    FOREIGN BONDPADCNU_m 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 34.100 BY 170.000 ;
    SYMMETRY X Y ;
    OBS
        LAYER metal4 ;
        RECT  -10.950 0.000 45.050 12.500 ;
        RECT  -10.950 15.500 45.050 28.500 ;
        RECT  -10.950 31.500 45.050 44.500 ;
        RECT  -10.950 0.000 7.050 60.000 ;
        RECT  10.050 0.000 24.050 60.000 ;
        RECT  27.050 0.000 45.050 60.000 ;
        RECT  5.550 67.000 28.550 82.000 ;
        RECT  5.550 89.000 28.550 104.000 ;
        RECT  5.550 111.000 28.550 126.000 ;
        RECT  5.550 133.000 28.550 148.000 ;
        RECT  5.550 47.500 14.740 170.000 ;
        RECT  19.360 47.500 28.550 170.000 ;
        RECT  5.550 155.000 28.550 170.000 ;
        LAYER metal5 ;
        RECT  -10.950 0.000 45.050 12.500 ;
        RECT  -10.950 15.500 45.050 28.500 ;
        RECT  -10.950 31.500 45.050 44.500 ;
        RECT  -10.950 0.000 7.050 60.000 ;
        RECT  10.050 0.000 24.050 60.000 ;
        RECT  27.050 0.000 45.050 60.000 ;
        RECT  5.550 67.000 28.550 82.000 ;
        RECT  5.550 89.000 28.550 104.000 ;
        RECT  5.550 111.000 28.550 126.000 ;
        RECT  5.550 133.000 28.550 148.000 ;
        RECT  5.550 47.500 14.740 170.000 ;
        RECT  19.360 47.500 28.550 170.000 ;
        RECT  5.550 155.000 28.550 170.000 ;
        LAYER metal6 ;
        RECT  -10.950 0.000 45.050 60.000 ;
        RECT  5.550 67.000 28.550 82.000 ;
        RECT  5.550 89.000 28.550 104.000 ;
        RECT  5.550 111.000 28.550 126.000 ;
        RECT  5.550 133.000 28.550 148.000 ;
        RECT  5.550 0.000 14.740 170.000 ;
        RECT  19.360 0.000 28.550 170.000 ;
        RECT  5.550 155.000 28.550 170.000 ;
    END
END BONDPADCNU_m

MACRO BONDPADCGU_m
    CLASS BLOCK ;
    FOREIGN BONDPADCGU_m 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 34.100 BY 66.000 ;
    SYMMETRY X Y ;
    OBS
        LAYER metal4 ;
        RECT  -10.950 0.000 45.050 12.500 ;
        RECT  -10.950 15.500 45.050 28.500 ;
        RECT  -10.950 31.500 45.050 44.500 ;
        RECT  -10.950 0.000 7.050 60.000 ;
        RECT  10.050 0.000 24.050 60.000 ;
        RECT  27.050 0.000 45.050 60.000 ;
        RECT  3.740 47.500 14.740 66.000 ;
        RECT  19.360 47.500 30.360 66.000 ;
        RECT  3.740 63.000 30.360 66.000 ;
        LAYER metal5 ;
        RECT  -10.950 0.000 45.050 12.500 ;
        RECT  -10.950 15.500 45.050 28.500 ;
        RECT  -10.950 31.500 45.050 44.500 ;
        RECT  -10.950 0.000 7.050 60.000 ;
        RECT  10.050 0.000 24.050 60.000 ;
        RECT  27.050 0.000 45.050 60.000 ;
        RECT  3.740 47.500 14.740 66.000 ;
        RECT  19.360 47.500 30.360 66.000 ;
        RECT  3.740 63.000 30.360 66.000 ;
        LAYER metal6 ;
        RECT  -10.950 0.000 45.050 60.000 ;
        RECT  3.740 0.000 14.740 66.000 ;
        RECT  19.360 0.000 30.360 66.000 ;
        RECT  3.740 63.000 30.360 66.000 ;
    END
END BONDPADCGU_m

END LIBRARY
