VERSION 5.5 ;
NAMESCASESENSITIVE ON ;





LAYER metal1  
    AntennaAreaRatio 400 ;
    AntennaCumAreaRatio 400 ;
    AntennaAreaFactor 1 ;  
END metal1

LAYER metal2
    AntennaAreaRatio 400 ;
    AntennaCumAreaRatio 400 ;
    AntennaAreaFactor 1 ;  
END metal2

LAYER metal3
    AntennaAreaRatio 400 ;
    AntennaCumAreaRatio 400 ;
    AntennaAreaFactor 1 ;  
END metal3

LAYER metal4  
    AntennaAreaRatio 400 ;
    AntennaCumAreaRatio 400 ;
    AntennaAreaFactor 1 ;  
END metal4

LAYER metal5  
    AntennaAreaRatio 400 ;
    AntennaCumAreaRatio 400 ;
    AntennaAreaFactor 1 ;  
END metal5

LAYER metal6
    AntennaAreaRatio 400 ;
    AntennaCumAreaRatio 400 ;
    AntennaAreaFactor 1 ;  
END metal6


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon Feb 12 16:30:26 CST 2007
#
#**********************************************************************




MACRO GNDIOC
  PIN GNDO
   AntennaPartialMetalArea                 2885.054000 LAYER metal5 ;
   AntennaPartialMetalArea                 2885.054000 LAYER metal6 ;
   AntennaDiffArea                          659.640000 LAYER metal5 ;
   AntennaDiffArea                          659.640000 LAYER metal6 ;
  END GNDO

END GNDIOC


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon Feb 12 16:30:32 CST 2007
#
#**********************************************************************




MACRO GNDIOD
  PIN GNDO
   AntennaPartialMetalArea                 2973.709400 LAYER metal5 ;
   AntennaPartialMetalArea                 2973.709400 LAYER metal6 ;
   AntennaDiffArea                          820.948000 LAYER metal5 ;
   AntennaDiffArea                          820.948000 LAYER metal6 ;
  END GNDO

END GNDIOD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon Jul 21 14:47:05 CST 2008
#
#**********************************************************************




MACRO VCC3IOC
  PIN VCC3O
   AntennaPartialMetalArea                 3069.194000 LAYER metal5 ;
   AntennaPartialMetalArea                 3069.194000 LAYER metal6 ;
   AntennaGateArea                          790.400000 LAYER metal5 ;
   AntennaGateArea                          790.400000 LAYER metal6 ;
   AntennaDiffArea                         2323.056800 LAYER metal5 ;
   AntennaDiffArea                         2323.056800 LAYER metal6 ;
   AntennaMaxAreaCAR                         18.252810 LAYER metal5 ; 
  END VCC3O

END VCC3IOC


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon Feb 12 16:30:21 CST 2007
#
#**********************************************************************




MACRO VCC3IOD
  PIN VCC3O
   AntennaPartialMetalArea                 3411.098000 LAYER metal5 ;
   AntennaPartialMetalArea                 3411.098000 LAYER metal6 ;
   AntennaGateArea                          969.200000 LAYER metal5 ;
   AntennaGateArea                          969.200000 LAYER metal6 ;
   AntennaDiffArea                         2231.695200 LAYER metal5 ;
   AntennaDiffArea                         2231.695200 LAYER metal6 ;
   AntennaMaxAreaCAR                         15.498401 LAYER metal5 ; 
  END VCC3O

END VCC3IOD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon Jul 21 14:45:29 CST 2008
#
#**********************************************************************




MACRO XMC
  PIN I
   AntennaPartialMetalArea                  130.204000 LAYER metal5 ;
   AntennaPartialMetalArea                  130.204000 LAYER metal6 ;
   AntennaDiffArea                         1639.282400 LAYER metal5 ;
   AntennaDiffArea                         1639.282400 LAYER metal6 ;
  END I

  PIN O
   AntennaPartialMetalArea                    6.775200 LAYER metal1 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaDiffArea                            2.430000 LAYER metal1 ;
   AntennaDiffArea                            2.430000 LAYER metal2 ;
   AntennaDiffArea                            2.430000 LAYER metal3 ;
  END O

  PIN PD
   AntennaPartialMetalArea                    5.366400 LAYER metal1 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.288000 LAYER metal1 ;
   AntennaGateArea                            0.288000 LAYER metal2 ;
   AntennaGateArea                            0.288000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          2.842567 LAYER metal1 ; 
  END PD

  PIN PU
   AntennaPartialMetalArea                    6.380000 LAYER metal1 ;
   AntennaPartialMetalArea                    2.963200 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.468000 LAYER metal1 ;
   AntennaGateArea                            0.576000 LAYER metal2 ;
   AntennaGateArea                            0.576000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          2.325921 LAYER metal1 ; 
  END PU

  PIN SMT
   AntennaPartialMetalArea                    4.905800 LAYER metal1 ;
   AntennaPartialMetalArea                    5.830400 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.288000 LAYER metal1 ;
   AntennaGateArea                            1.308000 LAYER metal2 ;
   AntennaGateArea                            1.308000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          2.842572 LAYER metal1 ; 
  END SMT

END XMC


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon Jul 21 14:50:08 CST 2008
#
#**********************************************************************




MACRO XMD
  PIN I
   AntennaPartialMetalArea                  170.760000 LAYER metal5 ;
   AntennaPartialMetalArea                  170.760000 LAYER metal6 ;
   AntennaDiffArea                         1639.259600 LAYER metal5 ;
   AntennaDiffArea                         1639.259600 LAYER metal6 ;
  END I

  PIN O
   AntennaPartialMetalArea                    5.796000 LAYER metal1 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaDiffArea                            2.430000 LAYER metal1 ;
   AntennaDiffArea                            2.430000 LAYER metal2 ;
   AntennaDiffArea                            2.430000 LAYER metal3 ;
  END O

  PIN PD
   AntennaPartialMetalArea                    4.346400 LAYER metal1 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.288000 LAYER metal1 ;
   AntennaGateArea                            0.288000 LAYER metal2 ;
   AntennaGateArea                            0.288000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          2.842633 LAYER metal1 ; 
  END PD

  PIN PU
   AntennaPartialMetalArea                    3.072800 LAYER metal1 ;
   AntennaPartialMetalArea                    5.295600 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.180000 LAYER metal1 ;
   AntennaGateArea                            0.576000 LAYER metal2 ;
   AntennaGateArea                            0.576000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          1.747789 LAYER metal1 ; 
  END PU

  PIN SMT
   AntennaPartialMetalArea                    4.353800 LAYER metal1 ;
   AntennaPartialMetalArea                    5.654000 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.288000 LAYER metal1 ;
   AntennaGateArea                            1.308000 LAYER metal2 ;
   AntennaGateArea                            1.308000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          2.842639 LAYER metal1 ; 
  END SMT

END XMD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon Jul 21 14:48:47 CST 2008
#
#**********************************************************************




MACRO YA2GSC
  PIN E
   AntennaPartialMetalArea                    6.672800 LAYER metal1 ;
   AntennaPartialMetalArea                    5.945200 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.450000 LAYER metal1 ;
   AntennaGateArea                            1.350000 LAYER metal2 ;
   AntennaGateArea                            1.350000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          1.525556 LAYER metal1 ; 
  END E

  PIN E2
   AntennaPartialMetalArea                    6.920000 LAYER metal1 ;
   AntennaPartialMetalArea                    9.033600 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.288000 LAYER metal1 ;
   AntennaGateArea                            1.138000 LAYER metal2 ;
   AntennaGateArea                            1.138000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          2.542622 LAYER metal1 ; 
  END E2

  PIN E4
   AntennaPartialMetalArea                    5.852000 LAYER metal1 ;
   AntennaPartialMetalArea                   14.588800 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.288000 LAYER metal1 ;
   AntennaGateArea                            1.138000 LAYER metal2 ;
   AntennaGateArea                            1.138000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          2.542556 LAYER metal1 ; 
  END E4

  PIN E8
   AntennaPartialMetalArea                    6.344000 LAYER metal1 ;
   AntennaPartialMetalArea                    8.137600 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.288000 LAYER metal1 ;
   AntennaGateArea                            1.138000 LAYER metal2 ;
   AntennaGateArea                            1.138000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          2.542622 LAYER metal1 ; 
  END E8

  PIN I
   AntennaPartialMetalArea                    5.076800 LAYER metal1 ;
   AntennaPartialMetalArea                    7.544000 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.450000 LAYER metal1 ;
   AntennaGateArea                            1.350000 LAYER metal2 ;
   AntennaGateArea                            1.350000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          1.525522 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                  130.204000 LAYER metal5 ;
   AntennaPartialMetalArea                  130.204000 LAYER metal6 ;
   AntennaDiffArea                         1644.142000 LAYER metal5 ;
   AntennaDiffArea                         1644.142000 LAYER metal6 ;
  END O

  PIN SR
   AntennaPartialMetalArea                    4.975200 LAYER metal1 ;
   AntennaPartialMetalArea                    7.121200 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.384000 LAYER metal1 ;
   AntennaGateArea                            1.744000 LAYER metal2 ;
   AntennaGateArea                            1.744000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          2.094450 LAYER metal1 ; 
  END SR

END YA2GSC


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon Jul 21 14:49:23 CST 2008
#
#**********************************************************************




MACRO YA2GSD
  PIN E
   AntennaPartialMetalArea                    4.409600 LAYER metal1 ;
   AntennaPartialMetalArea                    7.880000 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            1.350000 LAYER metal2 ;
   AntennaGateArea                            1.350000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          5.121963 LAYER metal2 ; 
  END E

  PIN E2
   AntennaPartialMetalArea                    5.640800 LAYER metal1 ;
   AntennaPartialMetalArea                    6.460400 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.288000 LAYER metal1 ;
   AntennaGateArea                            1.138000 LAYER metal2 ;
   AntennaGateArea                            1.138000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          2.542589 LAYER metal1 ; 
  END E2

  PIN E4
   AntennaPartialMetalArea                    4.592000 LAYER metal1 ;
   AntennaPartialMetalArea                    6.872000 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.288000 LAYER metal1 ;
   AntennaGateArea                            1.138000 LAYER metal2 ;
   AntennaGateArea                            1.138000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          2.542556 LAYER metal1 ; 
  END E4

  PIN E8
   AntennaPartialMetalArea                    5.048000 LAYER metal1 ;
   AntennaPartialMetalArea                    5.312400 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.288000 LAYER metal1 ;
   AntennaGateArea                            1.138000 LAYER metal2 ;
   AntennaGateArea                            1.138000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          2.542622 LAYER metal1 ; 
  END E8

  PIN I
   AntennaPartialMetalArea                    4.724000 LAYER metal1 ;
   AntennaPartialMetalArea                    8.630400 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.450000 LAYER metal1 ;
   AntennaGateArea                            1.350000 LAYER metal2 ;
   AntennaGateArea                            1.350000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          1.525522 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                  170.760000 LAYER metal5 ;
   AntennaPartialMetalArea                  170.760000 LAYER metal6 ;
   AntennaDiffArea                         1644.142000 LAYER metal5 ;
   AntennaDiffArea                         1644.142000 LAYER metal6 ;
  END O

  PIN SR
   AntennaPartialMetalArea                    5.484800 LAYER metal1 ;
   AntennaPartialMetalArea                    9.067200 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.384000 LAYER metal1 ;
   AntennaGateArea                            1.744000 LAYER metal2 ;
   AntennaGateArea                            1.744000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          2.094467 LAYER metal1 ; 
  END SR

END YA2GSD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon Jul 21 14:47:36 CST 2008
#
#**********************************************************************




MACRO ZMA2GSC
  PIN E
   AntennaPartialMetalArea                    4.227200 LAYER metal1 ;
   AntennaPartialMetalArea                   11.702000 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            1.638000 LAYER metal2 ;
   AntennaGateArea                            1.638000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                         15.196322 LAYER metal2 ; 
  END E

  PIN E2
   AntennaPartialMetalArea                    6.920000 LAYER metal1 ;
   AntennaPartialMetalArea                    9.033600 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.288000 LAYER metal1 ;
   AntennaGateArea                            1.138000 LAYER metal2 ;
   AntennaGateArea                            1.138000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          2.542622 LAYER metal1 ; 
  END E2

  PIN E4
   AntennaPartialMetalArea                    5.852000 LAYER metal1 ;
   AntennaPartialMetalArea                   14.684000 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.288000 LAYER metal1 ;
   AntennaGateArea                            1.138000 LAYER metal2 ;
   AntennaGateArea                            1.138000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          2.542556 LAYER metal1 ; 
  END E4

  PIN E8
   AntennaPartialMetalArea                    6.344000 LAYER metal1 ;
   AntennaPartialMetalArea                    8.137600 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.288000 LAYER metal1 ;
   AntennaGateArea                            1.138000 LAYER metal2 ;
   AntennaGateArea                            1.138000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          2.542622 LAYER metal1 ; 
  END E8

  PIN I
   AntennaPartialMetalArea                    5.076800 LAYER metal1 ;
   AntennaPartialMetalArea                    7.544000 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.450000 LAYER metal1 ;
   AntennaGateArea                            1.350000 LAYER metal2 ;
   AntennaGateArea                            1.350000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          1.525522 LAYER metal1 ; 
  END I

  PIN IO
   AntennaPartialMetalArea                  130.204000 LAYER metal5 ;
   AntennaPartialMetalArea                  130.204000 LAYER metal6 ;
   AntennaDiffArea                         1639.282400 LAYER metal5 ;
   AntennaDiffArea                         1639.282400 LAYER metal6 ;
  END IO

  PIN O
   AntennaPartialMetalArea                    6.775200 LAYER metal1 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaDiffArea                            2.430000 LAYER metal1 ;
   AntennaDiffArea                            2.430000 LAYER metal2 ;
   AntennaDiffArea                            2.430000 LAYER metal3 ;
  END O

  PIN PD
   AntennaPartialMetalArea                    5.366400 LAYER metal1 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.288000 LAYER metal1 ;
   AntennaGateArea                            0.288000 LAYER metal2 ;
   AntennaGateArea                            0.288000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          2.842567 LAYER metal1 ; 
  END PD

  PIN PU
   AntennaPartialMetalArea                    3.663200 LAYER metal1 ;
   AntennaPartialMetalArea                    5.250800 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.180000 LAYER metal1 ;
   AntennaGateArea                            0.576000 LAYER metal2 ;
   AntennaGateArea                            0.576000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          1.405589 LAYER metal1 ; 
  END PU

  PIN SMT
   AntennaPartialMetalArea                    4.905800 LAYER metal1 ;
   AntennaPartialMetalArea                    5.830400 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.288000 LAYER metal1 ;
   AntennaGateArea                            1.308000 LAYER metal2 ;
   AntennaGateArea                            1.308000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          2.842572 LAYER metal1 ; 
  END SMT

  PIN SR
   AntennaPartialMetalArea                    4.975200 LAYER metal1 ;
   AntennaPartialMetalArea                    7.121200 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.384000 LAYER metal1 ;
   AntennaGateArea                            1.744000 LAYER metal2 ;
   AntennaGateArea                            1.744000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          2.094450 LAYER metal1 ; 
  END SR

END ZMA2GSC


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon Jul 21 14:45:47 CST 2008
#
#**********************************************************************




MACRO ZMA2GSD
  PIN E
   AntennaPartialMetalArea                    4.409600 LAYER metal1 ;
   AntennaPartialMetalArea                   13.312000 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            1.638000 LAYER metal2 ;
   AntennaGateArea                            1.638000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                         15.196316 LAYER metal2 ; 
  END E

  PIN E2
   AntennaPartialMetalArea                    5.640800 LAYER metal1 ;
   AntennaPartialMetalArea                    6.460400 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.288000 LAYER metal1 ;
   AntennaGateArea                            1.138000 LAYER metal2 ;
   AntennaGateArea                            1.138000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          2.542589 LAYER metal1 ; 
  END E2

  PIN E4
   AntennaPartialMetalArea                    4.592000 LAYER metal1 ;
   AntennaPartialMetalArea                    6.872000 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.288000 LAYER metal1 ;
   AntennaGateArea                            1.138000 LAYER metal2 ;
   AntennaGateArea                            1.138000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          2.542556 LAYER metal1 ; 
  END E4

  PIN E8
   AntennaPartialMetalArea                    5.048000 LAYER metal1 ;
   AntennaPartialMetalArea                    5.312400 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.288000 LAYER metal1 ;
   AntennaGateArea                            1.138000 LAYER metal2 ;
   AntennaGateArea                            1.138000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          2.542622 LAYER metal1 ; 
  END E8

  PIN I
   AntennaPartialMetalArea                    4.724000 LAYER metal1 ;
   AntennaPartialMetalArea                    8.630400 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.450000 LAYER metal1 ;
   AntennaGateArea                            1.350000 LAYER metal2 ;
   AntennaGateArea                            1.350000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          1.525522 LAYER metal1 ; 
  END I

  PIN IO
   AntennaPartialMetalArea                  170.760000 LAYER metal5 ;
   AntennaPartialMetalArea                  170.760000 LAYER metal6 ;
   AntennaDiffArea                         1639.259600 LAYER metal5 ;
   AntennaDiffArea                         1639.259600 LAYER metal6 ;
  END IO

  PIN O
   AntennaPartialMetalArea                    5.796000 LAYER metal1 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaDiffArea                            2.430000 LAYER metal1 ;
   AntennaDiffArea                            2.430000 LAYER metal2 ;
   AntennaDiffArea                            2.430000 LAYER metal3 ;
  END O

  PIN PD
   AntennaPartialMetalArea                    4.346400 LAYER metal1 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.288000 LAYER metal1 ;
   AntennaGateArea                            0.288000 LAYER metal2 ;
   AntennaGateArea                            0.288000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          2.842633 LAYER metal1 ; 
  END PD

  PIN PU
   AntennaPartialMetalArea                    3.111200 LAYER metal1 ;
   AntennaPartialMetalArea                    5.250800 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.180000 LAYER metal1 ;
   AntennaGateArea                            0.576000 LAYER metal2 ;
   AntennaGateArea                            0.576000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          1.405556 LAYER metal1 ; 
  END PU

  PIN SMT
   AntennaPartialMetalArea                    4.353800 LAYER metal1 ;
   AntennaPartialMetalArea                    5.654000 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.288000 LAYER metal1 ;
   AntennaGateArea                            1.308000 LAYER metal2 ;
   AntennaGateArea                            1.308000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          2.842639 LAYER metal1 ; 
  END SMT

  PIN SR
   AntennaPartialMetalArea                    5.484800 LAYER metal1 ;
   AntennaPartialMetalArea                    9.067200 LAYER metal2 ;
   AntennaPartialMetalArea                    1.692000 LAYER metal3 ;
   AntennaGateArea                            0.384000 LAYER metal1 ;
   AntennaGateArea                            1.744000 LAYER metal2 ;
   AntennaGateArea                            1.744000 LAYER metal3 ;
   AntennaDiffArea                            0.490000 LAYER metal1 ;
   AntennaDiffArea                            0.490000 LAYER metal2 ;
   AntennaDiffArea                            0.490000 LAYER metal3 ;
   AntennaMaxAreaCAR                          2.094467 LAYER metal1 ; 
  END SR

END ZMA2GSD

END LIBRARY
